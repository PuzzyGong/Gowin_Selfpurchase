//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18C
//Created Time: Tue Oct 25 12:42:16 2022

module ROM_varies (dout, clk, oce, ce, reset, ad);

output [0:0] dout;
input clk;
input oce;
input ce;
input reset;
input [14:0] ad;

wire lut_f_0;
wire lut_f_1;
wire [30:0] prom_inst_0_dout_w;
wire [0:0] prom_inst_0_dout;
wire [30:0] prom_inst_1_dout_w;
wire [0:0] prom_inst_1_dout;
wire dff_q_0;

LUT2 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[14])
);
defparam lut_inst_0.INIT = 4'h2;
LUT2 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[14])
);
defparam lut_inst_1.INIT = 4'h8;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],prom_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hE3F8FCFFE3F8FCFFE000FCFFF7FCFCFFFFFFF8FFFFFFFCFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_01 = 256'hE3F8C03FE3F8F07FE3F8FC7FE000FC7FE3F8FCFFE3F80003E3F89CFFE3F8FCFF;
defparam prom_inst_0.INIT_RAM_02 = 256'hE3F8FCF7E3F8FCE7E3F8FCCFE3F8FCCFE000FC9FE3F8DC1FE3F8CC3FE3F8C43F;
defparam prom_inst_0.INIT_RAM_03 = 256'hFFFFFFFFFFFCFEFFE3F8FCFFE3F8FCFFE000FCFFE3F8FCFFE3F8FCF9E3F8FCFB;
defparam prom_inst_0.INIT_RAM_04 = 256'hFE7E7E7FFE7E7E7FFC007E7FFE7F7E7FFFFFFC7FFFFFFF7FFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_05 = 256'hFE7E701FFE7E7C3FFE7E7E3FFE7E7E3FFE7E7E3FFE7E4003FE7E667FFE7E7E7F;
defparam prom_inst_0.INIT_RAM_06 = 256'hCE7F3E7BCE7F3E73FE7E3E67FE7E7E67FE7E7E4FFE7E4E0FFE7E461FFE7E621F;
defparam prom_inst_0.INIT_RAM_07 = 256'hFFFFFFFFFFFFFF7FFFFFF27FC07FE67F807FCE7FCE7FCE7FCE7F9E7FCE7F1E7D;
defparam prom_inst_0.INIT_RAM_08 = 256'hFFCFEE7F800FFE7FCFCFFE7FFFCFFE7FFF8FFC7FFFEFFF7FFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_09 = 256'hF38E4663F3CE4663F3FE4663F3FE4663E0004663FBCFC663FFCFC663FFCF8003;
defparam prom_inst_0.INIT_RAM_0A = 256'hF3E67E7FF3CE7673F3CE6263F3CE4463F3CE4663F3CE4663F3CE4663F3CE4663;
defparam prom_inst_0.INIT_RAM_0B = 256'hFFFFFFFFFFFFC77FE7FF9E7FC7FE7E7FE3F8FE7FF1F1FE7FFCF3FE7FFF27FE7F;
defparam prom_inst_0.INIT_RAM_0C = 256'hFFFF3FFFE0000007F3FE7FFFFFFE7FFFFFFE3FFFFFFF9FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0D = 256'hFF9F3DFFFFFE7FFFFF9CE37FFF38027FFE71E63FF0E3CF1FF8F79FCFFFFE1FFF;
defparam prom_inst_0.INIT_RAM_0E = 256'h80000001E7FE7FFFFFFE7FFFFFEC7FEFF3CF43C7F1C00387F0E7CF3FFC739CFF;
defparam prom_inst_0.INIT_RAM_0F = 256'hFFFFFFFFFFFE7FFFFFFE7FFFFFFE7FFFFFFE7FFFFFFE7FFFFFFE7FFFFFFE7FFF;
defparam prom_inst_0.INIT_RAM_10 = 256'hFE3FFC7FFE3FFC7FFE3FFC7FFC00007FFF7FFF7FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_11 = 256'hFE3FFC7FFE00007FFE3FFC7FFE3FFC7FFE3FFC7FFE3FFC7FFE00007FFE3FFC7F;
defparam prom_inst_0.INIT_RAM_12 = 256'hFF33C43FFE73C63FFCF3C71FF8F3C79FE1F3C7EFF3F3C7FFFFE387FFFFFFFF7F;
defparam prom_inst_0.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFC0000003E3F3C7FFFFE3C7FFFFC3C67FFF93C47F;
defparam prom_inst_0.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFF800001FFC7FFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_15 = 256'hFFFE7FFFFFFE7FFF80000001E7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_16 = 256'hF1FE7F9FF8FE7F3FFC7E7E3FFE7E7C7FFF3E78FFFFDE70FFFFEE79FFFFFE7FFF;
defparam prom_inst_0.INIT_RAM_17 = 256'hFFFFFFFFFFFF9FFFFFFE1FFFFFFE07FFFFFE39F9E7FE7FF3E3FE7FE7E3FE7FCF;
defparam prom_inst_0.INIT_RAM_18 = 256'hFFCFEE7F800FFE7FCFCFFE7FFFCFFE7FFF8FFC7FFFEFFF7FFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_19 = 256'hF38E4663F3CE4663F3FE4663F3FE4663E0004663FBCFC663FFCFC663FFCF8003;
defparam prom_inst_0.INIT_RAM_1A = 256'hF3E67E7FF3CE7673F3CE6263F3CE4463F3CE4663F3CE4663F3CE4663F3CE4663;
defparam prom_inst_0.INIT_RAM_1B = 256'hFFFFFFFFFFFFC77FE7FF9E7FC7FE7E7FE3F8FE7FF1F1FE7FFCF3FE7FFF27FE7F;
defparam prom_inst_0.INIT_RAM_1C = 256'hFFFF3FFFE0000007F3FE7FFFFFFE7FFFFFFE3FFFFFFF9FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1D = 256'hFF9F3DFFFFFE7FFFFF9CE37FFF38027FFE71E63FF0E3CF1FF8F79FCFFFFE1FFF;
defparam prom_inst_0.INIT_RAM_1E = 256'h80000001E7FE7FFFFFFE7FFFFFEC7FEFF3CF43C7F1C00387F0E7CF3FFC739CFF;
defparam prom_inst_0.INIT_RAM_1F = 256'hFFFFFFFFFFFE7FFFFFFE7FFFFFFE7FFFFFFE7FFFFFFE7FFFFFFE7FFFFFFE7FFF;
defparam prom_inst_0.INIT_RAM_20 = 256'hF3FE7C7FF3FE7C7FE0007E3FFBFF7F3FFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_21 = 256'hF3FE7E7FF3FE7E7FF3FE7C01F3FE7F7FF3FE7FFFF3FE7FFFF3FE7FFFF3FE7EFF;
defparam prom_inst_0.INIT_RAM_22 = 256'hFCE0F67FFE61EE7FFFFBDE7FFFFFFE7FF3FE7E7FF3FE7E7FF0007E7FF3FE7E7F;
defparam prom_inst_0.INIT_RAM_23 = 256'hFFFFFFFFFFFFF7FFCFFFEFFFC7FF9E7FC7FF3C3FE3FE3C7FE1FC787FF9F8F27F;
defparam prom_inst_0.INIT_RAM_24 = 256'hE3CE3F9FE3FE3F9FE3FE3F9FE3FE001FE3FE7FDFF3FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_25 = 256'hE3CFF9FFE3CFF9FFE3CFF1DFE3CE399FE3CE001FE3CE3F9FE3CE3F9FE38E3F9F;
defparam prom_inst_0.INIT_RAM_26 = 256'hE3CE7E7FE3CE7CFFE3CC7CFFE3CC7CFFE3CC78FFE3CC79FFE3C80003E3CCF9FF;
defparam prom_inst_0.INIT_RAM_27 = 256'hFFFFFFFFF9FFDFFBF0FF1FF3E03F07EFE3FE3B9FE3FE7F1FE3FE7F3FE3FE7E7F;
defparam prom_inst_0.INIT_RAM_28 = 256'hFFF3FF1FC000011FF3F3FF8FFFF3FFE7FFE3FFFFFFF3FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_29 = 256'hF8000F3FF8F3CF3FF8F3CE01F8F3CF3FF8F3CFFFF0000FFFFDF3EFFFFFF3FFBF;
defparam prom_inst_0.INIT_RAM_2A = 256'hF3F3E73FF1F3CF3FF0F39F3FFC733F3FFF027F3FFFE0FF3FFFF1EF3FF8F1CF3F;
defparam prom_inst_0.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFE0007FFFC0000FF3BFFFE3F1FFF3F9E3FFF3FCCFFFF3FA1F;
defparam prom_inst_0.INIT_RAM_2C = 256'hFFFF3FFFE0000007F3FE7FFFFFFE7FFFFFFE3FFFFFFF9FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2D = 256'hFF9F3DFFFFFE7FFFFF9CE37FFF38027FFE71E63FF0E3CF1FF8F79FCFFFFE1FFF;
defparam prom_inst_0.INIT_RAM_2E = 256'h80000001E7FE7FFFFFFE7FFFFFEC7FEFF3CF43C7F1C00387F0E7CF3FFC739CFF;
defparam prom_inst_0.INIT_RAM_2F = 256'hFFFFFFFFFFFE7FFFFFFE7FFFFFFE7FFFFFFE7FFFFFFE7FFFFFFE7FFFFFFE7FFF;
defparam prom_inst_0.INIT_RAM_30 = 256'hFF8FFDFFC0000003E3FC7FFFFFFC7FFFFFFE3FFFFFFF9FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_31 = 256'hF90FE78FF9C3878FF9FBCF8FF9FFFF8FF000000FFBF7E7FFFFE7E3FFFFCFF3FF;
defparam prom_inst_0.INIT_RAM_32 = 256'hF9E7E78FF9E7E78FF9E7E78FF9E7E78FF9C0070FF9E7F48FF93FF98FF91FF38F;
defparam prom_inst_0.INIT_RAM_33 = 256'hFFFFFFFFFCFFFFCFF87FFF8FF81FFF8FF9F7E78FF9E7E78FF9E0078FF9E7E78F;
defparam prom_inst_0.INIT_RAM_34 = 256'hFF9FF9FFFF9FF9FFFF9FF9FFFF9FF9FFFF0001FFFF9FFDFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_35 = 256'hFFFFFFFFFFDFF9FFFF9FF9FFFF8001FFFF9FF9FFFF9FF9FFFF9FF9FFFF9FF9FF;
defparam prom_inst_0.INIT_RAM_36 = 256'hF3F1CFCFF3F1CFCFF3F1CFCFF3F1CFCFF3F1CFCFF3F1CFCFE001800FF3F9EFEF;
defparam prom_inst_0.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFEFFBF1FFCFF3F1CFCFF3F1CFCFF001C00FF3F1CFCFF3F1CFCF;
defparam prom_inst_0.INIT_RAM_38 = 256'hFFFBCFFFFFF3C7FFFFE7C7FFFFC7E3FFFF87F3FFFFEFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_39 = 256'hFE7FFC7FFE7FFC7FFE7FFC7FFE7FFC7FFE7FFC7FFE7FFC7FFC00007FFE79FF7F;
defparam prom_inst_0.INIT_RAM_3A = 256'hF1BCF1DFFE7C71FFFFFC79FFFFFF1F7FFE7FDC7FFE00007FFE7FFC7FFE7FFC7F;
defparam prom_inst_0.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFF8003FFFF0001FFFF9FF1E3E7BFF1C3E3BFF1C7E3BFF1CF;
defparam prom_inst_0.INIT_RAM_3C = 256'hFFE7C93FFFE7991FFFC7399FFFC639CFFF8FF1FFFFEFF9FFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3D = 256'hF8E6F9E7F8F4398FF9F5191FF9F1803FF9F1E07FF9F3F8FF80000003E7F269FF;
defparam prom_inst_0.INIT_RAM_3E = 256'hFF1FCE1FFE1FCF3FFE1F9E7FFE4F9E7FFC4F0003FCEFBCFFFCEFF8FFFCE77DF3;
defparam prom_inst_0.INIT_RAM_3F = 256'hFFFFFFFFFFFF8FFFE7FE3FE183FCFF8FE0F27E7FF8E638FFFC0F03FFFE1FC1FF;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[30:0],prom_inst_1_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 1;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hFF8FFDFFC0000003E3FC7FFFFFFC7FFFFFFE3FFFFFFF9FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_01 = 256'hF90FE78FF9C3878FF9FBCF8FF9FFFF8FF000000FFBF7E7FFFFE7E3FFFFCFF3FF;
defparam prom_inst_1.INIT_RAM_02 = 256'hF9E7E78FF9E7E78FF9E7E78FF9E7E78FF9C0070FF9E7F48FF93FF98FF91FF38F;
defparam prom_inst_1.INIT_RAM_03 = 256'hFFFFFFFFFCFFFFCFF87FFF8FF81FFF8FF9F7E78FF9E7E78FF9E0078FF9E7E78F;
defparam prom_inst_1.INIT_RAM_04 = 256'hFF9FF9FFFF9FF9FFFF9FF9FFFF9FF9FFFF0001FFFF9FFDFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_05 = 256'hFFFFFFFFFFDFF9FFFF9FF9FFFF8001FFFF9FF9FFFF9FF9FFFF9FF9FFFF9FF9FF;
defparam prom_inst_1.INIT_RAM_06 = 256'hF3F1CFCFF3F1CFCFF3F1CFCFF3F1CFCFF3F1CFCFF3F1CFCFE001800FF3F9EFEF;
defparam prom_inst_1.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFEFFBF1FFCFF3F1CFCFF3F1CFCFF001C00FF3F1CFCFF3F1CFCF;
defparam prom_inst_1.INIT_RAM_08 = 256'hFFFBCFFFFFF3C7FFFFE7C7FFFFC7E3FFFF87F3FFFFEFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_09 = 256'hFE7FFC7FFE7FFC7FFE7FFC7FFE7FFC7FFE7FFC7FFE7FFC7FFC00007FFE79FF7F;
defparam prom_inst_1.INIT_RAM_0A = 256'hF1BCF1DFFE7C71FFFFFC79FFFFFF1F7FFE7FDC7FFE00007FFE7FFC7FFE7FFC7F;
defparam prom_inst_1.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFF8003FFFF0001FFFF9FF1E3E7BFF1C3E3BFF1C7E3BFF1CF;
defparam prom_inst_1.INIT_RAM_0C = 256'hFFCCFE7FFFE8FC7FFFE1FC7FFFF1FCFFFFE1F8FFFFFBFCFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0D = 256'hFF3E7837E63C722783FF660FE0FFCE1FF87F9E1FFE7F3F1FFF3E3F3FFF9C7E3F;
defparam prom_inst_1.INIT_RAM_0E = 256'hFF3F3E3FFF3E3E3FFF3E7E3FFF3E7E3FFF3E7E3FFF3E7E3FFF3E7E39FF3E7E33;
defparam prom_inst_1.INIT_RAM_0F = 256'hFFBFFFBFFF3FF83FFF3FF63FFF3FCE3FFF3F8E3FFF3F9E3FFF3F3E3FFF3F3E3F;
defparam prom_inst_1.INIT_RAM_10 = 256'hF9FE7F1FF9FE7F1FF9FE7F1FF9FE7F1FF000001FFBFFFF9FFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_11 = 256'hF9FE7F1FF9FE7F1FF9FE7F1FF9FE7F1FF800001FF9FE7F1FF9FE7F1FF9FE7F1F;
defparam prom_inst_1.INIT_RAM_12 = 256'hF9FE7FCFF9FE7F9FF9FE7F9FF9FE7F9FF9FE7F9FF800001FF9FE7F9FF9FE7F9F;
defparam prom_inst_1.INIT_RAM_13 = 256'hFFFFFFFFFCFFFFF9F8FFFFFBF83E7FF3F80E7FE7F9FE7FE7F9FE7FCFF9FE7FCF;
defparam prom_inst_1.INIT_RAM_14 = 256'hF000007FF9FCFE7FFFF8FFFFFFFC7FFFFFFE7FFFFFFF3FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_15 = 256'hF80000FFF8FFFCFFF8FFFCFFF8FFFCFFF8FFFCFFF8FFFCFFF8FFFCFFF8FFFCFF;
defparam prom_inst_1.INIT_RAM_16 = 256'hFFFFFF3FFFFFFE3FFFFFFE7FFFFFFE7FFFFFFE7FFFFFFC7FF8FFFC7FF8FFFCFF;
defparam prom_inst_1.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFF9FFFFFFF3FFFFFFE7FFFFFFCFFFFFFFCFFFFFFF9FFFFFFF1F;
defparam prom_inst_1.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_20 = 256'hEFF1C7E7FFF3C7E7FFF3C007FFE3EFFFFFC3FFFFFFF7FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_21 = 256'hE7E38667E7E70667E7C74667C7F64667C7FCC667C7FCC667C7F9C467C001C767;
defparam prom_inst_1.INIT_RAM_22 = 256'hE7FEFD3FE4F06627E4024667E67CC667E73DC667E799C667E7F3C667E7F3C667;
defparam prom_inst_1.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFDF8FFFFF3F03F9FE7F39F9FCFE3FF8FDFE7FFC79FE7FFF33F;
defparam prom_inst_1.INIT_RAM_24 = 256'hFCF9FCFFF9FFFFFFC1FFFFFFE000000FF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_25 = 256'hFFF9F8FFFFF9FC7FFFF9FE7FFFF9FF9FFFF9CFFFFFF9C7FFFF79C7FFFEF1F3FF;
defparam prom_inst_1.INIT_RAM_26 = 256'hFFE63FFFFFF87FFFFFFCFFFFFFFCFFFFC0000003E7F8FFFFFFF8F9FFFFF9F9FF;
defparam prom_inst_1.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFC3F3FFFF1FE1FFF8FFF0FFF3FFF07FC7FFFC3F8FFFFF0F1FFF;
defparam prom_inst_1.INIT_RAM_28 = 256'hFFF9C7FFFFFC8FFFFFFE1FFFFFFF1FFFFFFE3FFFFFFF3FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_29 = 256'hE3FE3FE78100009FE01FFE3FFC3FFC7FFF0FF8FFFFC7F1FFFFE7E3FFFFF3C7FF;
defparam prom_inst_1.INIT_RAM_2A = 256'hFE1E3E7FFF9E3F7FFFFE3FFFF800001FFCFE3FFFFFFE3FFFFFFE3FFFFFFE3FF1;
defparam prom_inst_1.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFC0000003E7F633FFFFE633FFFFCE31FFFF8E31FFFF9E38FF;
defparam prom_inst_1.INIT_RAM_2C = 256'hFFDF3FE7FF9E0007FF9F39EFFF1FF9FF80007CFFEFFFFE7FFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2D = 256'hE739F0E7E739F20FE639E7CFE7B9E79FE7F9C01FE7F9EF3FC001DE33E7DF9F63;
defparam prom_inst_1.INIT_RAM_2E = 256'hFE1DCF9FE799CF99E799CF83E739C00FE739FF9FE7391F3FE7398E7FE739C0F3;
defparam prom_inst_1.INIT_RAM_2F = 256'hFFFFFFFFDFFF1FFFCFFE7F9FCFF9EF9FC7F3C01FE3E7CF9FF1CFCF9FFC8FCF9F;
defparam prom_inst_1.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_0 (
  .O(dout[0]),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_1_dout[0]),
  .S0(dff_q_0)
);
endmodule //ROM_varies
