//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18C
//Created Time: Wed Oct 26 16:44:38 2022

module ROM_character (dout, clk, oce, ce, reset, ad);

output [0:0] dout;
input clk;
input oce;
input ce;
input reset;
input [14:0] ad;

wire lut_f_0;
wire lut_f_1;
wire [30:0] prom_inst_0_dout_w;
wire [0:0] prom_inst_0_dout;
wire [30:0] prom_inst_1_dout_w;
wire [0:0] prom_inst_1_dout;
wire dff_q_0;

LUT2 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[14])
);
defparam lut_inst_0.INIT = 4'h2;
LUT2 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[14])
);
defparam lut_inst_1.INIT = 4'h8;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],prom_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0C = 256'hFFFFE7E7FFFF8381FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0D = 256'hFFFFFE7FFFFFFC3FFFFFFD3FFFFFF91FFFFFFB9FFFFFF38FFFFFF3CFFFFFE7CF;
defparam prom_inst_0.INIT_RAM_0E = 256'hFFFFFE7FFFFFFE7FFFFFFE7FFFFFFE7FFFFFFE7FFFFFFE7FFFFFF00FFFFFFE7F;
defparam prom_inst_0.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF81FFFFFFE7FFFFFFE7FFFFFFE7F;
defparam prom_inst_0.INIT_RAM_10 = 256'hFFFF1FFFFFFF1FFFFFFF1FFFFFFF1FFFFFFE1FFFFFFF9FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_11 = 256'hFFFF187FFFFF07FFFFF81FFFFF871FFFF87F1FFFC3FF1FFFF3FF1FFFFFFF1FFF;
defparam prom_inst_0.INIT_RAM_12 = 256'hEFFF1FFFEFFF1FFFEFFF1FFFEFFF1FFFFFFF1FFFFFFF1FFFFFFF1FF1FFFF1F87;
defparam prom_inst_0.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFC0003FFF80001FFFC7FF1FFFE7FF1FFFE7FF1FFF;
defparam prom_inst_0.INIT_RAM_14 = 256'hFFFE7FFFFFFE7FFFF000000FF8FE7FFFFFFC7FFFFFFF7FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_15 = 256'hFF3FFCFFFF3FFCFFFF3FFCFFFE0000FFFF3FFFFFFFFFFFFFFE00007FFF3E7FFF;
defparam prom_inst_0.INIT_RAM_16 = 256'hFE0000FFFF7FFEFFC0000003E3F3CFFFFFE7CFFFFFC7E7FFFF27FCFFFF0000FF;
defparam prom_inst_0.INIT_RAM_17 = 256'hFFFFFFFFFF3FFCFFFF3FFCFFFF0000FFFF3FFCFFFF3FFCFFFF3FFCFFFF3FFCFF;
defparam prom_inst_0.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1C = 256'hE3C7E7E7F81F8381FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1D = 256'hE3FFFE7FE7FFFC3FC7FFFD3FC7E3F91FC7E3FB9FC7F3F38FC7F3F3CFE7E3E7CF;
defparam prom_inst_0.INIT_RAM_1E = 256'hDFE7FE7FDFCFFE7FFF9FFE7FFF3FFE7FFE7FFE7FFCFFFE7FF9FFF00FF1FFFE7F;
defparam prom_inst_0.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC001F81FC001FE7FCFF3FE7FCFF3FE7F;
defparam prom_inst_0.INIT_RAM_20 = 256'hFFFF3FFFFFFE3FFFFFFE3FFFC0000003F3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_21 = 256'hFE3FFC7FFE3FFC7FFE3FFC7FFE3FFC7FFC00007FFE7F9F7FFFFF9FFFFFFF3FFF;
defparam prom_inst_0.INIT_RAM_22 = 256'hFE3FFC7FFE3FFC7FFE3FFC7FFE3FFC7FFE00007FFE3FFC7FFE3FFC7FFE3FFC7F;
defparam prom_inst_0.INIT_RAM_23 = 256'hFFFFFFFFFF3FFE7FFE3FFC7FFE3FFC7FFE00007FFE3FFC7FFE3FFC7FFE3FFC7F;
defparam prom_inst_0.INIT_RAM_24 = 256'hFFFE7FFFFFFE7FFFC0000003E3FE7FFFFFFC7FFFFFFE7FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_25 = 256'hFE7E7FFFFE7E7E7FFE00007FFE7E7E7FFE7E7E7FFE7E7E7FFC00007FFEFE7FFF;
defparam prom_inst_0.INIT_RAM_26 = 256'hFE7E7FFFFE7E7FFFFE7E7FFF80000001E67E7FFFFE7E7FFFFE7E7FFFFC00001F;
defparam prom_inst_0.INIT_RAM_27 = 256'hFFFFFFFFFFFFBFFFFFFE1FFFFFFE03FFFFFE7FFFFF7E7FFFFE7E7FFFFE00001F;
defparam prom_inst_0.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2C = 256'hE3C7E7E7F81F8381FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2D = 256'hE3FFFE7FE7FFFC3FC7FFFD3FC7E3F91FC7E3FB9FC7F3F38FC7F3F3CFE7E3E7CF;
defparam prom_inst_0.INIT_RAM_2E = 256'hDFE7FE7FDFCFFE7FFF9FFE7FFF3FFE7FFE7FFE7FFCFFFE7FF9FFF00FF1FFFE7F;
defparam prom_inst_0.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC001F81FC001FE7FCFF3FE7FCFF3FE7F;
defparam prom_inst_0.INIT_RAM_30 = 256'hFF3E7C7FFEFE78FFFDFE7FFFE1FE7FFFE000000FF3FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_31 = 256'hFFFC7FFBF07E7FF78001FFCFFFF83F9FFFFE4F9FFFFE673FFFFE783FFE007C7F;
defparam prom_inst_0.INIT_RAM_32 = 256'hFC00003FFCFE7E3FFCFE7E3FFCFE7E3FFCFE7E3FFCFE7E3FF800003FFCFE7FBF;
defparam prom_inst_0.INIT_RAM_33 = 256'hFFFFFFFFE7FFFFEFE7FFF807E3C00007F01E7FFFFC7E7FFFFF3E7FFFFEFE7E3F;
defparam prom_inst_0.INIT_RAM_34 = 256'hFFE7E3FFE000000FF9E7E3FFFFE7E3FFFFC7E3FFFFF7F3FFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_35 = 256'hFE7E7E7FFC00007FFEFE7FFFFFFE7FFF80000001C7E7E3FFFFE7E3FFFFE7E3FF;
defparam prom_inst_0.INIT_RAM_36 = 256'hFE00007FFE7E7E7FFE7E7E7FFE7E7E7FFE7E7E7FFE00007FFE7E7E7FFE7E7E7F;
defparam prom_inst_0.INIT_RAM_37 = 256'hFFFFFFFFF3FFFFF3F1FFFF8FF0FFFE3FF87FFC7FFF1FF1FFFFE3C3FFFE7FE67F;
defparam prom_inst_0.INIT_RAM_38 = 256'hFBFF9A7FFFFF9E7FFFF01E7FF00FFE3FF07FFF1FFBFFFFDFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_39 = 256'hF8D99E7FC3D99ECFE7D99CCFFFD99DC7FFD99DC7FFC19DF3FC1D9BF9F0FF9BFF;
defparam prom_inst_0.INIT_RAM_3A = 256'hFC79E78FFE79C78FFF39CF81FF39CF1FFF39CF3FFF99CF3FFF998F7FFE198E7F;
defparam prom_inst_0.INIT_RAM_3B = 256'hFFFFFFFFFFFFFF7FFFF9FEFFC7F0FD8F83E1F98FE1C9F38FF8B9F38FFCF9E78F;
defparam prom_inst_0.INIT_RAM_3C = 256'hE3C7E7E7F81F8381FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3D = 256'hE3FFFE7FE7FFFC3FC7FFFD3FC7E3F91FC7E3FB9FC7F3F38FC7F3F3CFE7E3E7CF;
defparam prom_inst_0.INIT_RAM_3E = 256'hDFE7FE7FDFCFFE7FFF9FFE7FFF3FFE7FFE7FFE7FFCFFFE7FF9FFF00FF1FFFE7F;
defparam prom_inst_0.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC001F81FC001FE7FCFF3FE7FCFF3FE7F;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[30:0],prom_inst_1_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 1;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hFF1FFE7FFC3FFE3FFC00063FFE7FFF1FFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_01 = 256'hE739DCDFC0000D8FE7FE1D87FFFC79C7FFF8FBF3FFF3FBFFFFE7F3FFFFCFFFFF;
defparam prom_inst_1.INIT_RAM_02 = 256'hF3E3E38FE3E7CF83E3C79F1FE3CF3F3FE38E3F3FE79C7E7FE71CFE7FE738FEFF;
defparam prom_inst_1.INIT_RAM_03 = 256'hFFFFFFFFFE7FF9FFF83FE38FF80F8F8FF1E73F8FF3FC7F8FF3F8FE9FF3F1F99F;
defparam prom_inst_1.INIT_RAM_04 = 256'hFFF3FFFFFFE3FE7FFFE3FE7FFFE3FE3FFFE3FF9FFFF3FFDFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_05 = 256'hFFF9FF3FFFF1FF3FFFF3FE01FFF3FF3FFFF3FFFFC00003FFE7F3FFFFFFF3FFFF;
defparam prom_inst_1.INIT_RAM_06 = 256'hF3FFE73FF1FFCF3FF8FF9F3FF8FF3F3FFC7E7F3FFF3CFF3FFF98FF3FFFE1FF3F;
defparam prom_inst_1.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFE000FFFFC0000FF3BFFFC3F1FFFFF9E3FFFFFCCFFBFFFA1F;
defparam prom_inst_1.INIT_RAM_08 = 256'hFFFE3FFFFFFE3FFFFFFE3FFFFFFE3FFFFFFC3FFFFFFFBFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_09 = 256'hFFF98FFFFFF99FFFFFFD1FFFFFFC1FFFFFFC1FFFFFFC1FFFFFFE1FFFFFFE1FFF;
defparam prom_inst_1.INIT_RAM_0A = 256'hFF0FF1FFFF8FF3FFFFC7E3FFFFE7C7FFFFE3C7FFFFF3CFFFFFF38FFFFFF98FFF;
defparam prom_inst_1.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFF9F3FFFFE781FFFF8FE0FFFF1FF87FFE7FFC3FFCFFFF1FF8FF;
defparam prom_inst_1.INIT_RAM_0C = 256'hF1FFE7E7F3FF8381FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0D = 256'hF1CFFE7FF1DFFC3FF19FFD3FF13FF91FF17FFB9FF07FF38FF0FFF3CFF0FFE7CF;
defparam prom_inst_1.INIT_RAM_0E = 256'hF1FFFE7FF1FFFE7F8001FE7FF1F9FE7FF1FBFE7FF1F3FE7FF1E7F00FF1EFFE7F;
defparam prom_inst_1.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF803FF81FF1FFFE7FF1FFFE7FF1FFFE7F;
defparam prom_inst_1.INIT_RAM_10 = 256'hFFFCFF9FC000001FE3F9FFDFFFF9FFFFFFF8FFFFFFFE7FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_11 = 256'hFCF8FF9F8000001FE4F8FF9FFCF8FF9FFCF8FF9FF800019FFEF8FF9FFFF8FF9F;
defparam prom_inst_1.INIT_RAM_12 = 256'hFF981FCFFE48CFCFF8E8C79FE1E0E79FF3F0F99FFCF0FF9FFC00019FFCF8FF9F;
defparam prom_inst_1.INIT_RAM_13 = 256'hFFFFFFFFFFFE7FFDF7FC7FFBE1FC0EF3C0F8FC37FC78F0E7FE38E3E7FF988FCF;
defparam prom_inst_1.INIT_RAM_14 = 256'hFFCFFCC7FFCFFCE7FFCFFCFFC0000CFFE7FFF8FFFFFFFEFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_15 = 256'hE7CF9CC7E7CF9CC7E7CF9CC7E7CF9CC7E7CF9CC7C0001CC7F7CFDCC7FFCFFCC7;
defparam prom_inst_1.INIT_RAM_16 = 256'hE04F9F3FE7CF9E7FE7CF9E67E7CF9E47E7CF9C47E7CF9CC7E7CF9CC7E7CF9CC7;
defparam prom_inst_1.INIT_RAM_17 = 256'hFFFFFFFFFFEFFFF9FFCFFFF3FFCFFFE7FFCFFFCFFFCFFF9FFBCFFF9FF1CFDF3F;
defparam prom_inst_1.INIT_RAM_18 = 256'hC000023FE5F3FE7FFCF3FC7FFC73FCFFFE23F8FFFFF3FEFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_19 = 256'hF9F3CF37F9F3CF27F8000F0FF9F3CF0FF9F3CE1FF0000F1FF9F3FF3FFFF3FF3F;
defparam prom_inst_1.INIT_RAM_1A = 256'hFE7FBF3F8000013FE67FFF3FFC73CF3FFE73CF3FF9F3CF3FF8000F3FF9F3CF3B;
defparam prom_inst_1.INIT_RAM_1B = 256'hFFFFFFFFFF3FFFBFFE1FFF3FFE07FF3FFE7CFF3FFE7CFF3FFE7C7F3FFE7E7F3F;
defparam prom_inst_1.INIT_RAM_1C = 256'hF1E7E7E7FC1F8381FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1D = 256'hF9FFFE7FF3FFFC3FE3FFFD3FE7FFF91FE7E3FB9FE7E3F38FE3E3F3CFE3E3E7CF;
defparam prom_inst_1.INIT_RAM_1E = 256'hC7E3FE7FC7E3FE7FC7FFFE7FC7FFFE7FC7FFFE7FE3FFFE7FF1FFF00FFC3FFE7F;
defparam prom_inst_1.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF81FF81FF1E7FE7FE7E3FE7FC7E3FE7F;
defparam prom_inst_1.INIT_RAM_20 = 256'hFFE3FE7FFFE3C003FFE7E7FFC0003FFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_21 = 256'hF3FDFE7FC000FE7FF3F9FE7FFFF9FE7FFFF1FE7FFFF1FE7FFFF3FE7FFFF3FE7F;
defparam prom_inst_1.INIT_RAM_22 = 256'hF9FFFFC3F1FFFF03F1FFFC3FF3FFE07FF3FF8E7FF3FFFE7FF3FFFE7FF3FFFE7F;
defparam prom_inst_1.INIT_RAM_23 = 256'hFFFFFFFFFF1FFFFFFE1FFFFFFC07FFFFF8F3FFFFF8FFFFFFF9FFFFFFF9FFFFF7;
defparam prom_inst_1.INIT_RAM_24 = 256'hC0000003E3FE7FFFFFFE7FFFFFFE7FFFFFFC7FFFFFFE7FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_25 = 256'hFF3FFC7FFF3FFC7FFF3FFC7FFF3FFC7FFE00007FFF7E7FFFFFFE7FFFFFFE7FFF;
defparam prom_inst_1.INIT_RAM_26 = 256'hEFF1C7FFFFF1CFFFFFF1CFFFFFF1CE7FFF31CC7FFF00007FFF3FFC7FFF3FFC7F;
defparam prom_inst_1.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFE3E003FF1FC3F3FC7FE7F1F9FFE7F1F3FFE7F1E3FFEFF1E7FF;
defparam prom_inst_1.INIT_RAM_28 = 256'hFFFE7FFFFFFE7FFFFFFE7FFFFFFE7FFFFFFC7FFFFFFF7FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_29 = 256'hF3FF1FFFF3FF3FFFF3FF3FFFF3FE3FFFF3FE3FFFE000000FF3FE7FFFFFFE7FFF;
defparam prom_inst_1.INIT_RAM_2A = 256'hF9FFF1FFF9FFE3FFF9FFE7FFF1FFC7FFF1FFCFFFF1FF8FFFF1FF9FFFF1FF1FFF;
defparam prom_inst_1.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFF9FF1FFFE7FE0FFF8FFC03FF3FFCF9FE7FF8FFFCFFF8FFF9FF;
defparam prom_inst_1.INIT_RAM_2C = 256'hE39FE7E7F03F8381FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2D = 256'hE391FE7FF031FC3FFFF3FD3FFFF3F91FFFE3FB9FFFE7F38FE7E7F3CFE3CFE7CF;
defparam prom_inst_1.INIT_RAM_2E = 256'hCFE3FE7FCFF3FE7F8FF3FE7F8FF1FE7F8FF1FE7FCFF1FE7FCFE1F00FC7C1FE7F;
defparam prom_inst_1.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF81FF81FF38FFE7FE7C7FE7FCFE3FE7F;
defparam prom_inst_1.INIT_RAM_30 = 256'hFE7FFFFFFE7FFFFF80000001C3FFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_31 = 256'hFE7E7F3FFE7E7F3FFE7E7F3FFE7E7F3FFE7C003FFE7E7FBFFE7FFFFFFE7FFFFF;
defparam prom_inst_1.INIT_RAM_32 = 256'hFE7FFF3FFE7E7F3FFE7E7F3FFE7E003FFE7E7F3FFE7E7F3FFE7E7F3FFE7E7F3F;
defparam prom_inst_1.INIT_RAM_33 = 256'hFFFFFFFFFF9FFFFFFF1FFFFFFE03FFFFFE39FFFFFE7FFFFFFE7FFFFFFE7FFFFF;
defparam prom_inst_1.INIT_RAM_34 = 256'hF8FFFF3FF800003FFDFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_35 = 256'hF8FFFF3FF8FFFF3FF8FFFF3FF8FFFF3FF8FFFF3FF8FFFF3FF8FFFF3FF8FFFF3F;
defparam prom_inst_1.INIT_RAM_36 = 256'hF800003FF8FFFF3FF8FFFF3FF8FFFF3FF8FFFF3FF8FFFF3FF8FFFF3FF8FFFF3F;
defparam prom_inst_1.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFCFFFF3FF8FFFF3FF8FFFF3F;
defparam prom_inst_1.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3C = 256'hE3C7E7E7F81F8381FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3D = 256'hE3FFFE7FE7FFFC3FC7FFFD3FC7E3F91FC7E3FB9FC7F3F38FC7F3F3CFE7E3E7CF;
defparam prom_inst_1.INIT_RAM_3E = 256'hDFE7FE7FDFCFFE7FFF9FFE7FFF3FFE7FFE7FFE7FFCFFFE7FF9FFF00FF1FFFE7F;
defparam prom_inst_1.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC001F81FC001FE7FCFF3FE7FCFF3FE7F;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_0 (
  .O(dout[0]),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_1_dout[0]),
  .S0(dff_q_0)
);
endmodule //ROM_character
