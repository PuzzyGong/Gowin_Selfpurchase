//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18C
//Created Time: Sat Oct 01 22:14:30 2022

module ROM_letter_show (dout, clk, oce, ce, reset, ad);

output [0:0] dout;
input clk;
input oce;
input ce;
input reset;
input [13:0] ad;

wire [30:0] prom_inst_0_dout_w;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_10 = 256'h000000000000300033F800000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_11 = 256'h0000044004783FC0044004783FC0044000000006000C00100006000C00100000;
defparam prom_inst_0.INIT_RAM_12 = 256'h00001E0021181EE003001CF0210800F0000000001E302108FFFC208818700000;
defparam prom_inst_0.INIT_RAM_13 = 256'h00000000000000000000000E0016001010002100270019702488230821F01E00;
defparam prom_inst_0.INIT_RAM_14 = 256'h00000000000007E01818200440020000000040022004181807E0000000000000;
defparam prom_inst_0.INIT_RAM_15 = 256'h00000100010001001FF001000100010000000240024001800FF0018002400240;
defparam prom_inst_0.INIT_RAM_16 = 256'h01000100010001000100010001000000000000000000000000007000B0008000;
defparam prom_inst_0.INIT_RAM_17 = 256'h0004001800600180060018006000000000000000000000000000300030000000;
defparam prom_inst_0.INIT_RAM_18 = 256'h00000000200020003FF820102010000000000FE010102008200810100FE00000;
defparam prom_inst_0.INIT_RAM_19 = 256'h00000E3011482088208820081830000000003070218822082408280830700000;
defparam prom_inst_0.INIT_RAM_1A = 256'h00000E08110820882088210819F80000000024003FF82410242004C007000000;
defparam prom_inst_0.INIT_RAM_1B = 256'h00000008003800C83F0800080038000000000E0011182088208811100FE00000;
defparam prom_inst_0.INIT_RAM_1C = 256'h00000FE0111022082208311000E0000000001C7022882108210822881C700000;
defparam prom_inst_0.INIT_RAM_1D = 256'h0000000000000000608080000000000000000000000030C030C0000000000000;
defparam prom_inst_0.INIT_RAM_1E = 256'h0000044004400440044004400440044000002008101008200440028001000000;
defparam prom_inst_0.INIT_RAM_1F = 256'h000000F001083608300800480070000000000100028004400820101020080000;
defparam prom_inst_0.INIT_RAM_20 = 256'h20003800270002E0023823C03C00200000000BE0141023E8242827C8183007C0;
defparam prom_inst_0.INIT_RAM_21 = 256'h000008381008200820082008183007C000000E0011702088208820883FF82008;
defparam prom_inst_0.INIT_RAM_22 = 256'h00001810200823E8208820883FF8200800000FE010102008200820083FF82008;
defparam prom_inst_0.INIT_RAM_23 = 256'h000002001E38220820082008183007C000000010000803E8008820883FF82008;
defparam prom_inst_0.INIT_RAM_24 = 256'h00000000200820083FF820082008000020083FF821080100010021083FF82008;
defparam prom_inst_0.INIT_RAM_25 = 256'h000020083818262801C020883FF820080000000800087FF8800880088000C000;
defparam prom_inst_0.INIT_RAM_26 = 256'h000020083FF800F83F0000F83FF820080000300020002000200020083FF82008;
defparam prom_inst_0.INIT_RAM_27 = 256'h00000FE0101020082008200810100FE000083FF81808070000C020303FF82008;
defparam prom_inst_0.INIT_RAM_28 = 256'h00004FE0501038082408240818100FE0000000F001080108010821083FF82008;
defparam prom_inst_0.INIT_RAM_29 = 256'h00001C38220821082108208838700000200030700C880388008820883FF82008;
defparam prom_inst_0.INIT_RAM_2A = 256'h00081FF820082000200020081FF8000800000018000820083FF8200800080018;
defparam prom_inst_0.INIT_RAM_2B = 256'h000003F83C08070000F807003C0803F80008003801C80E003800078800780008;
defparam prom_inst_0.INIT_RAM_2C = 256'h00000008003820C83F0020C800380008200830182C68038003802C6830182008;
defparam prom_inst_0.INIT_RAM_2D = 256'h00004002400240027FFE00000000000000001808203820C82108260838082010;
defparam prom_inst_0.INIT_RAM_2E = 256'h0000000000007FFE40024002400200000000C0003800060001C00030000C0000;
defparam prom_inst_0.INIT_RAM_2F = 256'h8000800080008000800080008000800000000004000200020002000400000000;
defparam prom_inst_0.INIT_RAM_30 = 256'h20003F0022802280228024801900000000000000000000000004000200020000;
defparam prom_inst_0.INIT_RAM_31 = 256'h0000110020802080208011000E00000000000E0011002080208011003FF80008;
defparam prom_inst_0.INIT_RAM_32 = 256'h0000130022802280228022801F00000020003FF810882080208011000E000000;
defparam prom_inst_0.INIT_RAM_33 = 256'h0000608093809480948094806B00000000180088208820883FF0208020800000;
defparam prom_inst_0.INIT_RAM_34 = 256'h00000000200020003F9820982080000020003F0020800080008021003FF82008;
defparam prom_inst_0.INIT_RAM_35 = 256'h0000208030802D80020024003FF82008000000007F98809880808000C0000000;
defparam prom_inst_0.INIT_RAM_36 = 256'h3F00008020803F80008020803F80208000000000200020003FF8200820080000;
defparam prom_inst_0.INIT_RAM_37 = 256'h00001F0020802080208020801F00000020003F0020800080008021003F802080;
defparam prom_inst_0.INIT_RAM_38 = 256'h8000FF80A0802080208011000E00000000000E00110020802080A100FF808080;
defparam prom_inst_0.INIT_RAM_39 = 256'h00001980248024802480248033000000000001800080208021003F8020802080;
defparam prom_inst_0.INIT_RAM_3A = 256'h20003F8010802000200020001F80008000000000208020801FE0008000800000;
defparam prom_inst_0.INIT_RAM_3B = 256'h00800F8030800C0003800C0030800F80008001800680080030000E8001800080;
defparam prom_inst_0.INIT_RAM_3C = 256'h008001800680180070008E80818080800000208031800E802E00318020800000;
defparam prom_inst_0.INIT_RAM_3D = 256'h400240023F7C0080000000000000000000003080218022802C80308021800000;
defparam prom_inst_0.INIT_RAM_3E = 256'h00000000000000803F7C400240020000000000000000FFFF0000000000000000;
defparam prom_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000040004000200020001000100060000;

endmodule //ROM_letter_show
