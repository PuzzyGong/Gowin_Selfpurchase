//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18C
//Created Time: Tue Oct 25 13:56:58 2022

module ROM_ascii (dout, clk, oce, ce, reset, ad);

output [0:0] dout;
input clk;
input oce;
input ce;
input reset;
input [15:0] ad;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire [30:0] prom_inst_0_dout_w;
wire [0:0] prom_inst_0_dout;
wire [30:0] prom_inst_1_dout_w;
wire [0:0] prom_inst_1_dout;
wire [30:0] prom_inst_2_dout_w;
wire [0:0] prom_inst_2_dout;
wire [30:0] prom_inst_3_dout_w;
wire [0:0] prom_inst_3_dout;
wire dff_q_0;
wire dff_q_1;
wire mux_o_0;
wire mux_o_1;

LUT3 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15])
);
defparam lut_inst_0.INIT = 8'h02;
LUT3 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15])
);
defparam lut_inst_1.INIT = 8'h08;
LUT3 lut_inst_2 (
  .F(lut_f_2),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15])
);
defparam lut_inst_2.INIT = 8'h20;
LUT3 lut_inst_3 (
  .F(lut_f_3),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15])
);
defparam lut_inst_3.INIT = 8'h80;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],prom_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[30:0],prom_inst_1_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 1;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_02 = 256'hFE7FFE7FFE7FFE7FFE7FFE3FFE3FFE3FFE3FFE7FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFE3FFC3FFC3FFE3FFFFFFFFFFFFFFE7FFE7FFE7FFE7FFE7F;
defparam prom_inst_1.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF7BFEF7FCE7F9CFF18FE31FC21FE73FFFFFFFFF;
defparam prom_inst_1.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_06 = 256'hF7EFF7CF800180018001E7CFE7CFE7CFE7CFE7CFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFBE7FBE7F3E7F3E7F3E7800180018001F3E7F3EFF7EFF7EF;
defparam prom_inst_1.INIT_RAM_08 = 256'hFE1FFE0FFE47FE47E267E267E667E667F24FF83FFE7FFE7FFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_09 = 256'hFFFFFE7FFE7FFE7FFC1FF267E663E663C663C663C67FE67FE27FF07FF87FFC3F;
defparam prom_inst_1.INIT_RAM_0A = 256'hFE99FE9CFC9CFD9CF99CFB9CF39CF399F7D9E7E3FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFC3F799F799E79DEF9CCF9CDF9C9F9CBF99BF993FD943C249;
defparam prom_inst_1.INIT_RAM_0C = 256'hFF87FF27FE67FE67FCE7FCE7FCE7FCE7FE47FE0FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFC707807330F978F8F878FA38F238F318F799F789E783C1C7;
defparam prom_inst_1.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFE7FFCFFFCFFFCFFFC3FFC3FFC3FFFFFFFF;
defparam prom_inst_1.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_10 = 256'hFE7FFE7FFE7FFE7FFC7FFCFFFCFFF9FFF9FFF3FFF3FFE7FFCFFF9FFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_11 = 256'hFFFF9FFFCFFFE7FFF3FFF3FFF9FFF9FFFCFFFCFFFC7FFE7FFE7FFE7FFE7FFE7F;
defparam prom_inst_1.INIT_RAM_12 = 256'hFE7FFE7FFE7FFE3FFE3FFF3FFF3FFF9FFF9FFFCFFFE7FFE7FFF3FFF9FFFFFFFF;
defparam prom_inst_1.INIT_RAM_13 = 256'hFFFFFFF9FFF3FFE7FFE7FFCFFF9FFF9FFF3FFF3FFE3FFE3FFE7FFE7FFE7FFE7F;
defparam prom_inst_1.INIT_RAM_14 = 256'hFC3FF00FC24186618E71FE7FFC7FFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFE3FFE7F8E718661C241F00FFC3F;
defparam prom_inst_1.INIT_RAM_16 = 256'hFE7FFE7FFE7FFE7FFE7FFE7FFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFE7FFE7FFE7FFE7FFE7FFE7F8001;
defparam prom_inst_1.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_19 = 256'hFFF3FFE7FFCFFFCFFFCFFFC3FFC3FFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8001;
defparam prom_inst_1.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFC3FFC3FFC3FFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1E = 256'hFEFFFCFFFDFFF9FFFBFFF3FFF3FFE7FFE7FFCFFFCFFF9FFF9FFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1F = 256'hFFFFFFFFFFFDFFF9FFFBFFF3FFF7FFE7FFEFFFCFFFDFFF9FFFBFFF3FFF7FFE7F;
defparam prom_inst_1.INIT_RAM_20 = 256'h8FF18FF1CFF3C7F3C7E3C7E3E7E7E3C7F18FFC3FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFC3FF18FE3C7E7E7C7E3C7E3C7F3CFF3CFF18FF18FF18FF1;
defparam prom_inst_1.INIT_RAM_22 = 256'hFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE07FE7FFEFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFE007FC3FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7F;
defparam prom_inst_1.INIT_RAM_24 = 256'hE3FFE7FFC7FFC7E3C7E3C7F3C7F3E7E3E3C7F81FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFC001C001CFF3CFF3DFE7DFCFFF9FFF3FFE7FFCFFF9FFF1FF;
defparam prom_inst_1.INIT_RAM_26 = 256'hF9FFF3FFE3FFE7FFE7E3E7E3E3E3E3E3F1E7FC1FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFF81FF1E7E7E3C7E3C7E3C7E3C7FFC7FFC7FFE3FFF1FFFC3F;
defparam prom_inst_1.INIT_RAM_28 = 256'hF1CFF1DFF19FF13FF17FF07FF0FFF0FFF1FFF3FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFF803FF1FFF1FFF1FFF1FFF1FF8001F1F9F1FBF1F3F1E7F1EF;
defparam prom_inst_1.INIT_RAM_2A = 256'hF3C7F817FFF7FFF7FFF7FFF7FFF7FFF7C007C007FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFF81FF1E7E3F3C7F3C7E3CFE3CFFFCFFFCFFFC7FFC7F7E7E7;
defparam prom_inst_1.INIT_RAM_2C = 256'hE391F031FFF3FFF3FFE3FFE7E7E7E3CFE39FF03FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFF81FF38FE7C7CFE3CFE3CFF38FF38FF18FF1CFF1CFE1C7C1;
defparam prom_inst_1.INIT_RAM_2E = 256'hFCFFF9FFF9FFFBFFF3FBF7FBE7F3EFE3C003C007FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFE3FFE1FFE1FFE1FFE3FFE3FFE3FFE3FFE7FFE7FFE7FFCFF;
defparam prom_inst_1.INIT_RAM_30 = 256'hF00FE787E7E3CFF3CFF3CFF3CFF3E7E3E3C7F81FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFF81FF3C7E7F3CFF3CFF9CFF9CFF9C7F1C3F3E1E7F0CFF81F;
defparam prom_inst_1.INIT_RAM_32 = 256'hC7F1CFF1CFF1CFF1C7F1C7F1E7F3E3E3F1C7FC1FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFE0FF8C7F1E3F3E7E7FFE7FFC7FFC7FFC60FC1C7C3E3C7F3;
defparam prom_inst_1.INIT_RAM_34 = 256'hFC3FFC3FFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFE3FFC3FFC3FFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3F;
defparam prom_inst_1.INIT_RAM_36 = 256'hFC3FFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_37 = 256'hFFFFFF3FFE7FFE7FFC3FFC3FFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3F;
defparam prom_inst_1.INIT_RAM_38 = 256'hFFE7FFCFFF9FFF3FFE7FFCFFF9FFF3FFE7FFCFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFCFFFE7FFF3FFF9FFFCFFFE7FFF3FFF9FFFCFFFE7FFF3FFF3;
defparam prom_inst_1.INIT_RAM_3A = 256'hFFFFFFFF8001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8001FFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3C = 256'hE7FFF3FFF9FFFCFFFE7FFF3FFF9FFFCFFFE7FFF3FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFF3FFE7FFCFFF9FFF3FFE7FFCFFF9FFF3FFE7FFCFFFCFFF;
defparam prom_inst_1.INIT_RAM_3E = 256'hE3FFC7FFC7E38FE18FF18FFBCFF3C7F7E3CFF81FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFE3FFC3FFC3FFE3FFFFFFFFFFF7FFF7FFF7FFE7FFC7FF8FF;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[30:0],prom_inst_2_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 1;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'hB399B399B331B333A27380F39FE7CFCFE79FF83FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFF83FE78FCFE79FE7BFF3E233C893D9999999B399B399B399;
defparam prom_inst_2.INIT_RAM_02 = 256'hF9CFF9DFF8DFF89FFC9FFCBFFC3FFC3FFE3FFE7FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFF03E0C7F1C7F3E7F3E7F3E3F7E3F7E3E7F007F3EFF1EFF1CF;
defparam prom_inst_2.INIT_RAM_04 = 256'hF1E3E7E3C7E3C7E3C7E3C7E3C7E3C7E3E3E3F800FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFF000E3E3C7E38FE38FE38FE38FE38FE3CFE3C7E3E3E3F803;
defparam prom_inst_2.INIT_RAM_06 = 256'hFFF1FFF1FFF1FFF1BFF39FE39FE7CFC7C78FD83FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFF83FE78FCFC7DFE39FE3BFF1FFF1FFF1FFF1FFF1FFF1FFF1;
defparam prom_inst_2.INIT_RAM_08 = 256'h8FE38FE38FE38FE3CFE3C7E3C7E3E3E3F1E3FC00FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFC00F0E3E3E3E7E3C7E3CFE38FE38FE38FE38FE38FE38FE3;
defparam prom_inst_2.INIT_RAM_0A = 256'hF3E3F3E3F3E3FFE3FFE39FE3DFE3CFE3C7E3C001FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFC001C7E39FE39FE3BFE3FFE3FFE3FFE3F3E3F3E3F3E3F003;
defparam prom_inst_2.INIT_RAM_0C = 256'hF3E3F7E3F7E3FFE3FFE3BFE3BFE39FE387E3C001FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFF80FFE3FFE3FFE3FFE3FFE3FFE3F7E3F7E3F7E3F3E3F003;
defparam prom_inst_2.INIT_RAM_0E = 256'hFFF9FFF1FFF1FFF1CFF3CFF3EFE7E7C7E38FEC3FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFF81FF38FC7E7C7E3C7F3C7F1C7F1C7F1C7F901F9FFF9FFF9;
defparam prom_inst_2.INIT_RAM_10 = 256'hC7E3C7E3C7E3C7E3C7E3C7E3C7E3C7E3C7E303C0FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFF03C0C7E3C7E3C7E3C7E3C7E3C7E3C7E3C7E3C7E3C7E3C003;
defparam prom_inst_2.INIT_RAM_12 = 256'hFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FE007FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFE007FE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7F;
defparam prom_inst_2.INIT_RAM_14 = 256'hF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FF001FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_15 = 256'hFF03FC71FCF1F9F1F9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FF;
defparam prom_inst_2.INIT_RAM_16 = 256'hFE03FF23FF63FE63FCE3F9E3FBE3F3E3E7E38180FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFF0380C7E3E7E3E3E3E3E3F1E3F1E3F9E3F8E3FCE3FC43FE03;
defparam prom_inst_2.INIT_RAM_18 = 256'hFFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FF81FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFC001CFE79FE7BFE7BFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7;
defparam prom_inst_2.INIT_RAM_1A = 256'hC9CBC9C3CBC3C3C3C3E3C3E3C7E3C7E3C7F307F0FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFF0330CF3BCF3BCE3BCE1BCE1BCE1BCC9BCC9BCC8BCD8BC9CB;
defparam prom_inst_2.INIT_RAM_1C = 256'hDE3BDE3BDF1BDF1BDF8BDF83DFC3DFC3DFE303E0FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFCFC0CFFBC7FBC7FBC3FBC3FBC1FBD1FBD8FBD8FBDC7BDC7B;
defparam prom_inst_2.INIT_RAM_1E = 256'h8FF18FF18FF18FF18FF3CFE3C7E7E7C7F38FF83FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFF83FF38FE7C7C7E7CFE38FF38FF18FF18FF18FF18FF18FF1;
defparam prom_inst_2.INIT_RAM_20 = 256'hC7E38FE38FE38FE38FE38FE38FE3C7E3E3E3F001FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFF80FFE3FFE3FFE3FFE3FFE3FFE3FFE3FFE3FFE3F803E3E3;
defparam prom_inst_2.INIT_RAM_22 = 256'h8FF18FF18FF18FF18FF1CFF3C7E3E7C7F38FF81FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_23 = 256'hFFFFC7FFC3FFB1FFF01FF1CFE1E7C0E3CCC38E118FF18FF18FF18FF18FF18FF1;
defparam prom_inst_2.INIT_RAM_24 = 256'hE3E7C7E7C7E7CFE7CFE7CFE7C7E7C7E7E3E7F801FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFF0781C7E7E7E7E3E7E3E7F3E7F1E7F9E7F8E7F8E7FCE7F807;
defparam prom_inst_2.INIT_RAM_26 = 256'hFF0FFFC3FFE3FFF1CFF1CFF1E7F3E7F3E1E7FC1FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFF83BE3C3E7E3CFF3CFF9CFF9CFF9CFFFC7FFE1FFF07FFC1F;
defparam prom_inst_2.INIT_RAM_28 = 256'hFE7FFE7FFE7FFE7FFE7FBE7D9E7D9E79CE71C003FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFF80FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7F;
defparam prom_inst_2.INIT_RAM_2A = 256'hCFE3CFE3CFE3CFE3CFE3CFE3CFE3CFE3CFE303C0FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFF81FF3C7E7E7EFE3CFE3CFE3CFE3CFE3CFE3CFE3CFE3CFE3;
defparam prom_inst_2.INIT_RAM_2C = 256'hFBCFF3CFF7C7F7C7E7E7E7E7EFE3EFE3CFE383C0FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFF7FFE7FFE3FFE3FFE3FFC3FFC1FFD1FFD9FF99FF98FFB8F;
defparam prom_inst_2.INIT_RAM_2E = 256'hEC63EC73CC73CC73DC73DC73DE71DE719E710820FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFBCFFBCFF3CFF1CFF1CFF187F187F187E1A7E0A7E827EC27;
defparam prom_inst_2.INIT_RAM_30 = 256'hFE3FFC3FFD1FF99FFB8FF3CFF7C7E7E7E7E78381FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFF03C1C7E3E7E7E3EFF3CFF1DFF99FF89FF83FFC3FFC7FFE7F;
defparam prom_inst_2.INIT_RAM_32 = 256'hFD1FF99FFB8FF38FF3CFF7C7E7E7EFE3CFE38380FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFF80FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE3FFC3FFC1F;
defparam prom_inst_2.INIT_RAM_34 = 256'hFC7FFCFFF8FFF9FFF3FFE3FBE7F3C7F3CFC78007FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFC001C7F3CFE3DFE79FC7FFCFFF8FFF9FFF1FFF3FFE3FFE7F;
defparam prom_inst_2.INIT_RAM_36 = 256'hFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FC03FFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_37 = 256'hFFFFFFFFC03FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3FFF3F;
defparam prom_inst_2.INIT_RAM_38 = 256'hFF3FFF3FFF3FFF9FFF9FFFCFFFCFFFCFFFE7FFE7FFF3FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_39 = 256'hFFFF9FFFCFFFCFFFE7FFE7FFE7FFF3FFF3FFF9FFF9FFFCFFFCFFFCFFFE7FFE7F;
defparam prom_inst_2.INIT_RAM_3A = 256'hFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFC03FFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3B = 256'hFFFFFFFFFC03FCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFFFCFF;
defparam prom_inst_2.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7EFF18FF81FFC3FFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3F = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[30:0],prom_inst_3_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 1;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFF1FFF87FFFFFFFF;
defparam prom_inst_3.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_02 = 256'hE7E3F3E7F81FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFF8607A1E323F1E7F1E7F1E7F1E7E3E7C7E41FE3FFE7F3E7E3;
defparam prom_inst_3.INIT_RAM_04 = 256'hC7C3E383F063FFE3FFE3FFE3FFE3FFE3FFE3FFE0FFE7FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFF833F3C3E7E3C7E3CFE3CFE3CFE38FE3CFE3CFE3CFE3CFE3;
defparam prom_inst_3.INIT_RAM_06 = 256'hE7C7F38FF83FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFF81FE78FEFE7DFE3DFF3FFF3FFF3FFF3FFF3FFF3E7E3E7E7;
defparam prom_inst_3.INIT_RAM_08 = 256'hC7E7C1CFC41FC7FFC7FFC7FFC7FFC7FFC7FFC1FFCFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFE41F81CFC3E7C7E3C7F3C7F3C7F3C7F3C7F3C7F3C7E3C7E3;
defparam prom_inst_3.INIT_RAM_0A = 256'hE7C7F38FF83FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFF83FE78FEFE7DFE7FFE3FFF3FFF3C003CFF3CFF3CFE3C7E7;
defparam prom_inst_3.INIT_RAM_0C = 256'hFF1FFF1FE001FF1FFF1FFF1F9F3F9F3F8E7FC0FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFF003FF1FFF1FFF1FFF1FFF1FFF1FFF1FFF1FFF1FFF1FFF1F;
defparam prom_inst_3.INIT_RAM_0E = 256'hF3E781CF8C1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0F = 256'hF00FE7E7CFF3CFF3CFF3C7F3E00FFC07FFE7FFE7FC0FF1CFF3E7E7E3E7E3E7E7;
defparam prom_inst_3.INIT_RAM_10 = 256'hE7C3E383F063FFE3FFE3FFE3FFE3FFE3FFE3FFE1FFE7FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFF8181C7E3C7E3C7E3C7E3C7E3C7E3C7E3C7E3C7E3E7E3E7E3;
defparam prom_inst_3.INIT_RAM_12 = 256'hFE7FFE7FFE07FE7FFFFFFFFFFFFFFC7FFC3FFC7FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFE007FE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7F;
defparam prom_inst_3.INIT_RAM_14 = 256'hE3FFE3FFE07FE7FFFFFFFFFFFFFFE3FFE3FFE3FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_15 = 256'hFE07F9E3F3E3F3FFF3FFE3FFE3FFE3FFE3FFE3FFE3FFE3FFE3FFE3FFE3FFE3FF;
defparam prom_inst_3.INIT_RAM_16 = 256'hF9E7F3E7C0E7FFE7FFE7FFE7FFE7FFE7FFE7FFE1FFEFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFF8381C7E7E3E7F3E7F1E7F9E7F8C7FC07FE27FE67FEE7FCE7;
defparam prom_inst_3.INIT_RAM_18 = 256'hFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE07FE7FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFE007FE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7F;
defparam prom_inst_3.INIT_RAM_1A = 256'h9C718C61C300FFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFF00209E719E719E719E719E719E719E719E719E719E719E71;
defparam prom_inst_3.INIT_RAM_1C = 256'hE7C3E381F067FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFF8181C7E3C7E3C7E3C7E3C7E3C7E3C7E3C7E3C7E3E7E3E7E3;
defparam prom_inst_3.INIT_RAM_1E = 256'hE7E7F3CFF81FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFF81FF3CFE7E7CFF3CFF38FF18FF18FF18FF18FF1CFF3C7E3;
defparam prom_inst_3.INIT_RAM_20 = 256'hC7C3E381F827FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_21 = 256'hFF81FFE3FFE3FFE3F823E383E7E3CFE3CFE38FE38FE38FE38FE38FE3CFE3CFE3;
defparam prom_inst_3.INIT_RAM_22 = 256'hE3E7E1CFEC1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_23 = 256'h81FFE7FFE7FFE7FFE41FE1C7E3E7E7F3E7F3E7F3E7F1E7F1E7F1E7F3E7F3E7E3;
defparam prom_inst_3.INIT_RAM_24 = 256'h8E0F8C81C39FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFF801FF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF8FFF0F;
defparam prom_inst_3.INIT_RAM_26 = 256'hE7E7E3CFE81FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFF037E7C7CFE7CFF3CFF3C7FFE1FFF83FFE0FFFC7EFE7EFE7;
defparam prom_inst_3.INIT_RAM_28 = 256'hFF1FFF1FE003FF1FFF3FFF3FFF3FFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFF07FE63FEF3FDF3FFF3FFF1FFF1FFF1FFF1FFF1FFF1FFF1F;
defparam prom_inst_3.INIT_RAM_2A = 256'hE7E3E7E3E1E0EFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFE40F81C7E3E7E7E3E7E3E7E3E7E3E7E3E7E3E7E3E7E3E7E3;
defparam prom_inst_3.INIT_RAM_2C = 256'hE7E7E7E78381FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFE7FFE7FFE3FFC3FFC3FFD1FF99FF99FFB8FF3CFF7CFF7C7;
defparam prom_inst_3.INIT_RAM_2E = 256'hDE739E710400FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFBCFFBCFF1CFF18FF187F187E027E427EC23EC73CC73DE73;
defparam prom_inst_3.INIT_RAM_30 = 256'hF38FE7C7C103FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFF81C1E3E7E3EFF3CFF99FF8BFFC3FFC7FFE3FFC3FF91FFB9F;
defparam prom_inst_3.INIT_RAM_32 = 256'hE7C7E7C78181FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_33 = 256'hFFC3FF83FF3FFF3FFE7FFE7FFE7FFC7FFC3FFD3FF93FF99FFB9FF39FF3CFF7CF;
defparam prom_inst_3.INIT_RAM_34 = 256'hF3F3E3E3E003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFE003E7E3CFC7CFCFDF8FFF1FFF3FFE3FFC7FFCFFF8FBF1F3;
defparam prom_inst_3.INIT_RAM_36 = 256'hFCFFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFFBFFF3FFC7FFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_37 = 256'hFFFFC7FFF3FFFBFFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFFCFFFE3F;
defparam prom_inst_3.INIT_RAM_38 = 256'hFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7F;
defparam prom_inst_3.INIT_RAM_39 = 256'hFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7FFE7F;
defparam prom_inst_3.INIT_RAM_3A = 256'hFF3FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFFDFFFCFFFE3FFFFFFFF;
defparam prom_inst_3.INIT_RAM_3B = 256'hFFFFFFE3FFCFFFDFFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF9FFF3FFCFF;
defparam prom_inst_3.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE1FFD8FFBC7DBE39FF1BFF87FFFF;
defparam prom_inst_3.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[15]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_1_dout[0]),
  .S0(dff_q_1)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(prom_inst_2_dout[0]),
  .I1(prom_inst_3_dout[0]),
  .S0(dff_q_1)
);
MUX2 mux_inst_2 (
  .O(dout[0]),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_0)
);
endmodule //ROM_ascii
