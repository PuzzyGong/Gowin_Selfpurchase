`include "../define.v"

//16 个 长度为 16 (总32) 的字符串
//从左向右写，否则会覆盖
module const_str
#(
    parameter                           L_W = `LETTER_PIXEL_WIDTH   
)
(
    output             [16 * (32 * 8) - 1 : 0] o_str                       
);

assign o_str = {{ 109'b0,      3'b001, 8'd000, 8'd135, "FPS_1:          "} ,
                { 109'b0,      3'b010, 8'd000, 8'd155, "FPS_2:          "} ,
                { 109'b0,      3'b100, 8'd000, 8'd175, "faces:          "} ,
                { 109'b0,      3'b011, 8'd100, 8'd135, " Aaa :          "} ,
                { 109'b0,      3'b101, 8'd100, 8'd155, " Bbb :          "} ,
                { 109'b0,      3'b110, 8'd100, 8'd175, " Ccc :          "} ,
                { 109'b0,      3'b111, 8'd000, 8'd000, "                "} ,
                { 109'b0,      3'b111, 8'd000, 8'd000, "                "} ,
                { 109'b0,      3'b111, 8'd000, 8'd000, "                "} ,
                { 109'b0,      3'b111, 8'd000, 8'd000, "                "} ,
                { 109'b0,      3'b111, 8'd000, 8'd000, "                "} ,
                { 109'b0,      3'b111, 8'd000, 8'd000, "                "} ,
                { 109'b0,      3'b111, 8'd000, 8'd000, "                "} ,
                { 109'b0,      3'b111, 8'd000, 8'd000, "                "} ,
                { 109'b0,      3'b111, 8'd000, 8'd000, "                "} ,
                { 109'b0,      3'b111, 8'd000, 8'd000, "                "}};
                                    
endmodule