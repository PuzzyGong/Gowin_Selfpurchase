//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18C
//Created Time: Tue Oct 25 20:51:08 2022

module ROM_picture (dout, clk, oce, ce, reset, ad);

output [0:0] dout;
input clk;
input oce;
input ce;
input reset;
input [16:0] ad;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire [30:0] prom_inst_0_dout_w;
wire [0:0] prom_inst_0_dout;
wire [30:0] prom_inst_1_dout_w;
wire [0:0] prom_inst_1_dout;
wire [30:0] prom_inst_2_dout_w;
wire [0:0] prom_inst_2_dout;
wire [30:0] prom_inst_3_dout_w;
wire [0:0] prom_inst_3_dout;
wire [30:0] prom_inst_4_dout_w;
wire [0:0] prom_inst_4_dout;
wire [30:0] prom_inst_5_dout_w;
wire [0:0] prom_inst_5_dout;
wire [30:0] prom_inst_6_dout_w;
wire [0:0] prom_inst_6_dout;
wire [30:0] prom_inst_7_dout_w;
wire [0:0] prom_inst_7_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_0.INIT = 16'h0002;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_1.INIT = 16'h0008;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_2.INIT = 16'h0020;
LUT4 lut_inst_3 (
  .F(lut_f_3),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_3.INIT = 16'h0080;
LUT4 lut_inst_4 (
  .F(lut_f_4),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_4.INIT = 16'h0200;
LUT4 lut_inst_5 (
  .F(lut_f_5),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_5.INIT = 16'h0800;
LUT4 lut_inst_6 (
  .F(lut_f_6),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_6.INIT = 16'h2000;
LUT4 lut_inst_7 (
  .F(lut_f_7),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_7.INIT = 16'h8000;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],prom_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_01 = 256'hFFFFFFFFFF07FFFFFFFFFFFFFE07FFFFFFFFFFFFFF07FFFFFFFFFFFFFF87FFFF;
defparam prom_inst_0.INIT_RAM_02 = 256'hFFFFFFFF3FE1FFFFFFFFFFFFFFC3FFFFFFFFFFFFFF83FFFFFFFFFFFFFF83FFFF;
defparam prom_inst_0.INIT_RAM_03 = 256'hFF000FE7FC007FFFFFC07FFFE008FFFFFFF1FFFF00F0FFFFFFFFFFFC07E1FFFF;
defparam prom_inst_0.INIT_RAM_04 = 256'hFF83FF0FFE1F8FFFFF03FF8FFE1F1FFFFE03F807FC1E3FFFFE000007FE043FFF;
defparam prom_inst_0.INIT_RAM_05 = 256'hFFF1FF1FF803FFFFFFE3FF1F801FFFFFFFC3FF1C001FFFFFFFC3FF0E3E1FE7FF;
defparam prom_inst_0.INIT_RAM_06 = 256'hFFFFF01FC187F01FFFE0001FFD8F800FFFE01F1FFF0001FFFFF1FF1FFF003FFF;
defparam prom_inst_0.INIT_RAM_07 = 256'hFFFFFFFF0FE1FFFFFFFFFFFE07C3FFFFFFFFFF3F03C3FFFFFFFFFF3F0187FE7F;
defparam prom_inst_0.INIT_RAM_08 = 256'hFFFFE0007FFC3FFFFFFFF807FFF87FFFFFFFFC3FFFF0FFFFFFFFFFFF3FE1FFFF;
defparam prom_inst_0.INIT_RAM_09 = 256'hFFFFE0FFFE3FE3FFFFFFC07FFE1F87FFFFFFC07FF81F0FFFFFFFC03C001E1FFF;
defparam prom_inst_0.INIT_RAM_0A = 256'hFFFFE0C07E3FFFFFFFFFE0FFFE3FFFFFFFFFE0FFFE3FFFFFFFFFE0FFFE3FF9FF;
defparam prom_inst_0.INIT_RAM_0B = 256'hFFFFF0FFFC3FFFFFFFFFF0FFFC3FFFFFFFFFF0FE003FFFFFFFFFF0E0023FFFFF;
defparam prom_inst_0.INIT_RAM_0C = 256'hFFFFF0FFFC3FFFFFFFFFF0FFFC3FFFFFFFFFF0FFFC3FFFFFFFFFF0FFFC3FFFFF;
defparam prom_inst_0.INIT_RAM_0D = 256'hFFFFF03FFE3FFFFFFFFFF01C003FFFFFFFFFF000003FFFFFFFFFF0C0FC3FFFFF;
defparam prom_inst_0.INIT_RAM_0E = 256'hFFFFF87FFFFFFFFFFFFFF87FFE7FFFFFFFFFF03FFE7FFFFFFFFFF03FFE3FFFFF;
defparam prom_inst_0.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFFFFFF;
defparam prom_inst_0.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_11 = 256'hFFFFFFE07FE0FFFFFFFFFFF07FF0FFFFFFFFFFF83FFCFFFFFFFFFFFF7FFFFFFF;
defparam prom_inst_0.INIT_RAM_12 = 256'hFFFFE3F0FFF07FFFFFFFFFF0FFE07FFFFFFFFFF0FFC0FFFFFFFFFFF07FC0FFFF;
defparam prom_inst_0.INIT_RAM_13 = 256'hFFFFE038FF1E1FFFFFFF80F8FFDE1FFFFFFF81F8FFFC3FFFFFFF83F8FFF83FFF;
defparam prom_inst_0.INIT_RAM_14 = 256'hFFFDFFF8F07FE3FFFFFDFFE0F83FC7FFFFFFFF80FC3F8FFFFFFFFC08FE1F0FFF;
defparam prom_inst_0.INIT_RAM_15 = 256'hFFFCFFF0E0F0007FFFFCFFF8E08078FFFFFCFFF8E00FF1FFFFFDFFF8F07FE3FF;
defparam prom_inst_0.INIT_RAM_16 = 256'hFFF80001FFFFFC7FFFF80001FFFFF07FFFF83FE0F3FF803FFFF87FF0F1FE003F;
defparam prom_inst_0.INIT_RAM_17 = 256'hFFFFFFFC7E1FE3FFFFFFFFFFFC0003FFFFFFC01FFE007FFFFFFE0007FF07FFFF;
defparam prom_inst_0.INIT_RAM_18 = 256'hFFFF83F0FE1FE3FFFFFF87F0FE1FE3FFFFFFCFE0FE1FE3FFFFFFFFF07E1FE3FF;
defparam prom_inst_0.INIT_RAM_19 = 256'hFFFFF838FE1FE3FFFFFFC078FE1FE3FFFFFF00F0FE1003FFFFFF01F0FE1003FF;
defparam prom_inst_0.INIT_RAM_1A = 256'hFFBFFFF8FE1823FFFFFFFFE0FE1FE3FFFFFFFF80FE1FE3FFFFFFFE08FE1FE3FF;
defparam prom_inst_0.INIT_RAM_1B = 256'hFF9FFFF8FE1FF1FFFF9FFFF8FE1FF1FFFF9FFFF8FE1E71FFFFBFFFF8FE1001FF;
defparam prom_inst_0.INIT_RAM_1C = 256'hFF07FFE0FE1EF87FFF0FFFF0FE1FF07FFF0FFFF0FE1FF0FFFF1FFFF8FE1FF0FF;
defparam prom_inst_0.INIT_RAM_1D = 256'hFFC0000FFF07FC7FFF000003FE07F87FFE000001FE03F87FFE01FFC1FE01F87F;
defparam prom_inst_0.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFC007FFF0FFE7F;
defparam prom_inst_0.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_20 = 256'hFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_21 = 256'hFFFFFF81FE07FFFFFFFFFF80FF07FFFFFFFFFFC07FC7FFFFFFFFFFF07FF7FFFF;
defparam prom_inst_0.INIT_RAM_22 = 256'hFFFF87FFFFC1FFFFFFFFFFCFFF83FFFFFFFFFF87FF03FFFFFFFFFF83FE03FFFF;
defparam prom_inst_0.INIT_RAM_23 = 256'hFFFFFF8000307FFFFFFFF0000070FFFFFFFF0001FFE1FFFFFFFF003FFFC1FFFF;
defparam prom_inst_0.INIT_RAM_24 = 256'hFFFFFFC1FFF81FFFFFFFFFC1FFFC1FFFFFFFFFC1FFFC3FFFFFFFFFE000787FFF;
defparam prom_inst_0.INIT_RAM_25 = 256'hFFFFFF0000E1C3FFFFFFC00001E087FFFFFF8001FFF087FFFFFFC021FFF00FFF;
defparam prom_inst_0.INIT_RAM_26 = 256'hFFFFE3E1FFF1FE3FFFFFFFE1FFF1FC7FFFFFFFE1FFF1F0FFFFFFFFE103E1E1FF;
defparam prom_inst_0.INIT_RAM_27 = 256'hFFFFFFE000F1FFFFFFFFF0000071FFFFFFFF80007FF1FFCFFFFF8001FFF1FF1F;
defparam prom_inst_0.INIT_RAM_28 = 256'hFFF00FE1FFF0FFFFFFFFFFE1FFF0FFFFFFFFFFE1FFF1FFFFFFFFFFE1F7F1FFFF;
defparam prom_inst_0.INIT_RAM_29 = 256'hFFFFFFFF0000FFFFFFE0C0000000FFFFFFC0000007F0FFFFFFE00001FFF0FFFF;
defparam prom_inst_0.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFFF8FFFFFFFFFFFFFFF0FFFF;
defparam prom_inst_0.INIT_RAM_2B = 256'hFFFF00FC0001FFFFFFFF80000001FFFFFFFFC000FFFFFFFFFFFFF03FFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2C = 256'hFFFFE0FFFF87FFFFFFFFC0FFFF87FFFFFFFFC0FFFF83FFFFFFFF00FFFC03FFFF;
defparam prom_inst_0.INIT_RAM_2D = 256'hFFFFF001FF8FFFFFFFFFF87FFF8FFFFFFFFFF07FFF87FFFFFFFFF0FFFF87FFFF;
defparam prom_inst_0.INIT_RAM_2E = 256'hFFFFFFFFFF9FFFFFFFFFFFFFFF9FFFFFFFFFF000000FFFFFFFFFE000000FFFFF;
defparam prom_inst_0.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFF;
defparam prom_inst_0.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_31 = 256'hFFFFC3F0FF83FFFFFFFFF3E07FC3FFFFFFFFFFF07FE3FFFFFFFFFFFC7FFFFFFF;
defparam prom_inst_0.INIT_RAM_32 = 256'hFFFFF071FFF07FFFFFFFE0F0FFE0FFFFFFFF80F0FFC1FFFFFFFF81F0FF81FFFF;
defparam prom_inst_0.INIT_RAM_33 = 256'hFF9FFFC1FFF80FFFFF9FFF01FFFC1FFFFF9FFE01FFFC3FFFFFFFFC31FFF83FFF;
defparam prom_inst_0.INIT_RAM_34 = 256'hFE07FFC3C1F0F87FFF0FFFE00FF0F1FFFF0FFFE03FF0C3FFFF9FFFE07FF087FF;
defparam prom_inst_0.INIT_RAM_35 = 256'hFFFE007FFFF8FFFFFFC0000FFFF8FFEFFF000007FFF8FF9FFE00FF03F870FE3F;
defparam prom_inst_0.INIT_RAM_36 = 256'hFFFFF8007FF8FFFFFFFFFE07FFF8FFFFFFFFFFFFFFF8FFFFFFFFFFFFFFF8FFFF;
defparam prom_inst_0.INIT_RAM_37 = 256'hFFFFF87FFF87FFFFFFFFF83FFC03FFFFFFFFF03F0003FFFFFFFFF00003FDFFFF;
defparam prom_inst_0.INIT_RAM_38 = 256'hFFFFFC7E0787FFFFFFFFFC7F0787FFFFFFFFFC7FE787FFFFFFFFF87FFF87FFFF;
defparam prom_inst_0.INIT_RAM_39 = 256'hFFFFFC7F0F87FFFFFFFFFC7F0F87FFFFFFFFFC7F0F87FFFFFFFFFC7E0F87FFFF;
defparam prom_inst_0.INIT_RAM_3A = 256'hFFFFFC3F8787FFFFFFFFFC3F8787FFFFFFFFFC3F8F87FFFFFFFFFC3F0F87FFFF;
defparam prom_inst_0.INIT_RAM_3B = 256'hFFFFFEFFC3C7FFFFFFFFFC7FC7C7FFFFFFFFFC7F87C7FFFFFFFFFC3F87C7FFFF;
defparam prom_inst_0.INIT_RAM_3C = 256'hFFFFFF03F0FFFFFFFFFFFFE1E1FFFFFFFFFFFFFCE1FFFFFFFFFFFFFFC3EFFFFF;
defparam prom_inst_0.INIT_RAM_3D = 256'hFFFFC03FFE1FFFFFFFFFE01FFC3FFFFFFFFFF00FF87FFFFFFFFFFC07F0FFFFFF;
defparam prom_inst_0.INIT_RAM_3E = 256'hFFFF87FFFFF87FFFFFFF83FFFFE1FFFFFFFF81FFFF83FFFFFFFF80FFFF0FFFFF;
defparam prom_inst_0.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFF9FFFFFFE1FFF;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[30:0],prom_inst_1_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 1;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_01 = 256'hFFFFFFFFFFE07FFFFFFFFFFFFFF87FFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_02 = 256'hFFFFFFFFFFF0FFFFFFFFFFFFFFF0FFFFFFFFFFFFFFE0FFFFFFFFFFFFFFE07FFF;
defparam prom_inst_1.INIT_RAM_03 = 256'hFFFFFFFFFFF0FFFFFFFFFFFFFFF0FFFFFFFFFFFFFFF0FFFFFFFFFFFFFFF0FFFF;
defparam prom_inst_1.INIT_RAM_04 = 256'hFFFF001FFC30FFFFFFFF807FFFF0FFFFFFFFC0FFFFF0FFFFFFFFF1FFFFF0FFFF;
defparam prom_inst_1.INIT_RAM_05 = 256'hFFFFE1F83FC003FFFFFFE1F83E001FFFFFFFC1C01C007FFFFFFF80001800FFFF;
defparam prom_inst_1.INIT_RAM_06 = 256'hFFFFF0F87FF03FFFFFFFF1F87FF07007FFFFE1F87FF00007FFFFE1F83FF0003F;
defparam prom_inst_1.INIT_RAM_07 = 256'hFFFFF0FC7FF80FFFFFFFF0FC7FF01FFFFFFFF0F87FF01FFFFFFFF0F87FF03FFF;
defparam prom_inst_1.INIT_RAM_08 = 256'hFFFFF8FC3C0887FFFFFFF8FC7C0087FFFFFFF8FC7E000FFFFFFFF0FC7FF80FFF;
defparam prom_inst_1.INIT_RAM_09 = 256'hFDFFF0FE3FF8F0FFFDFFF0FC3FF8E1FFFFFFF8FC3C78C1FFFFFFF8FC3C18C3FF;
defparam prom_inst_1.INIT_RAM_0A = 256'hF8FFF0FF1FF8FE3FFCFFF0FE1FF8FC3FFCFFF0FE1FF8F87FFCFFF0FE1FF8F0FF;
defparam prom_inst_1.INIT_RAM_0B = 256'hF00803FFC3F87FF3F87F81FF87F87FC7F87FE1FF8FF87F8FF8FFE1FF0FF8FF1F;
defparam prom_inst_1.INIT_RAM_0C = 256'hFF807FFFFC783FFFF8001FFFF8F83FFFF00007FFF1F87FFFF00003FFE3F87FFF;
defparam prom_inst_1.INIT_RAM_0D = 256'hFFFFFFFFFFF87FFFFFFFFFFFFFF83FFFFFFFFFFFFFF83FFFFFFFFFFFFF383FFF;
defparam prom_inst_1.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFC7FFF;
defparam prom_inst_1.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_11 = 256'hFFFF8003FFFFFFFFFFFFC01FFFFFFFFFFFFFE07FFFFFFFFFFFFFF8FFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_12 = 256'hFFFFFFFF801FFFFFFFFFFFF801FFFFFFFFFFFF000FFFFFFFFFFFC000FFFFFFFF;
defparam prom_inst_1.INIT_RAM_13 = 256'hFFFFFFFE07FFFFFFFFFFFFFC0FFFFFFFFFFFFFFC0F803FFFFFFFFFFF0000FFFF;
defparam prom_inst_1.INIT_RAM_14 = 256'hFFFFF03FF87FFFFFFFFFF83FF0FFFFFFFFFFFC7FE1FFFFFFFFFFFFFF83FFFFFF;
defparam prom_inst_1.INIT_RAM_15 = 256'hFFFFFF81FF80FFFFFFFFFE07FF87FFFFFFFFFC0FFF0FFFFFFFFFF81FFE3FFFFF;
defparam prom_inst_1.INIT_RAM_16 = 256'hFFFFFFFE1FFCFFFFFFFFFFFC3FC07FFFFFFFFFF070007FFFFFFFFFE00000FFFF;
defparam prom_inst_1.INIT_RAM_17 = 256'hFFFFE07FF83FFFFFFFFFF83FE0FFFFFFFFFFFE3FC3FFFFFFFFFFFFFF07FFFFFF;
defparam prom_inst_1.INIT_RAM_18 = 256'hFFFF83FC00003FFFFFFF838000007FFFFFFFC000FF03FFFFFFFFC0FFFE1FFFFF;
defparam prom_inst_1.INIT_RAM_19 = 256'hFFFFFFFE1FFFFFFFFFFFFFFE1FFC3FFFFFFFCFFF0F801FFFFFFF87FFC0001FFF;
defparam prom_inst_1.INIT_RAM_1A = 256'hFFFFFE7E1FFDFFFFFFFFFFFE1FFFFFFFFFFFFFFE1FFFFFFFFFFFFFFE1FFFFFFF;
defparam prom_inst_1.INIT_RAM_1B = 256'hFFFC03FE1FFC1FFFFFFE01FE1FFC3FFFFFFF00FE1FFC7FFFFFFFC07E1FFCFFFF;
defparam prom_inst_1.INIT_RAM_1C = 256'hFFF83FFE1FFF03FFFFF81FFE1FFF07FFFFF80FFE1FFE07FFFFFC07FE1FFE0FFF;
defparam prom_inst_1.INIT_RAM_1D = 256'hFFFFFFFE00FFFFFFFFFFFFFE087FFFFFFFFFFFFE1FFFC7FFFFFCFFFE1FFF87FF;
defparam prom_inst_1.INIT_RAM_1E = 256'hFFFFFFFF07FFFFFFFFFFFFFF07FFFFFFFFFFFFFE03FFFFFFFFFFFFFE01FFFFFF;
defparam prom_inst_1.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFF;
defparam prom_inst_1.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_22 = 256'hFFFFF03FFFF07FFFFFFFF01FFFF07FFFFFFFF80FFFFC7FFFFFFFFE07FFFF7FFF;
defparam prom_inst_1.INIT_RAM_23 = 256'hFFFFFFFFFFFC3FFFFFFFFFFFFFFC3FFFFFFFF1FFFFF87FFFFFFFF07FFFF07FFF;
defparam prom_inst_1.INIT_RAM_24 = 256'hFFFF8003FC1F0FFFFFFC003FFF1F0FFFFFF803FFFFFE1FFFFFFE3FFFFFFE1FFF;
defparam prom_inst_1.INIT_RAM_25 = 256'hFFFFFF07FF07E1FFFFFFFF07FE0FC3FFFFFFFF800C0FC7FFFFFFF800081F87FF;
defparam prom_inst_1.INIT_RAM_26 = 256'hFFFF83E3FFF0003FFFFFE1C3FFE0003FFFFFFF87FFC3F87FFFFFFF07FF87F0FF;
defparam prom_inst_1.INIT_RAM_27 = 256'hFFFC00387FFE3FFFFFFC0FF8FFFC7FFFFFFE07F1FFF8FC3FFFFF07E1FFF8E03F;
defparam prom_inst_1.INIT_RAM_28 = 256'hFFFFF0E00FE003FFFFFFF87007838FFFFFFC7E400F1F0FFFFFFC38003FFF1FFF;
defparam prom_inst_1.INIT_RAM_29 = 256'hFFFFF8F0FFFFE1FFFFFFF8E1FFFF81FFFFFFF8C1FFFE01FFFFFFF0C18FF801FF;
defparam prom_inst_1.INIT_RAM_2A = 256'hF9FFFC7C1FC3FFFFFFFFF87C3F8FFFFFFFFFF8F87E3FFFFFFFFFF8F07FFFF3FF;
defparam prom_inst_1.INIT_RAM_2B = 256'hF9FFFC7FC3FF00FFF9FFFC7F87FE07FFF9FFFC7F0FF81FFFF9FFFC7E1FF0FFFF;
defparam prom_inst_1.INIT_RAM_2C = 256'hE01FE0FFFF1FFCFFF07FF0FFFC3FF07FF0FFF8FFF07FE01FF0FFF87FE1FFC01F;
defparam prom_inst_1.INIT_RAM_2D = 256'hFFE03FFFFFFFFFFFFE0007FFFFFFFFFFF80001FFFFF3FFFFE00001FFFFCFFFFF;
defparam prom_inst_1.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[30:0],prom_inst_2_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 1;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0A = 256'hFFFFFFFFFFFFF000000FFFFFFFFFFFFFFFFFFFFFFFFFFF8001FFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0B = 256'hFFFFFFFFFFFC000000003FFFFFFFFFFFFFFFFFFFFFFF80000001FFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0C = 256'hFFFFFFFFFFC00000000003FFFFFFFFFFFFFFFFFFFFF0000000000FFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0D = 256'hFFFFFFFFFE0000000000007FFFFFFFFFFFFFFFFFFF800000000001FFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0E = 256'hFFFFFFFFF00000000000000FFFFFFFFFFFFFFFFFFC0000000000003FFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0F = 256'hFFFFFFFFC000000000000003FFFFFFFFFFFFFFFFE000000000000007FFFFFFFF;
defparam prom_inst_2.INIT_RAM_10 = 256'hFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF8000000000000001FFFFFFFF;
defparam prom_inst_2.INIT_RAM_11 = 256'hFFFFFFFC00000000000000003FFFFFFFFFFFFFFE00000000000000007FFFFFFF;
defparam prom_inst_2.INIT_RAM_12 = 256'hFFFFFFF800000000000000001FFFFFFFFFFFFFF800000000000000001FFFFFFF;
defparam prom_inst_2.INIT_RAM_13 = 256'hFFFFFFE0000000000000000007FFFFFFFFFFFFF000000000000000000FFFFFFF;
defparam prom_inst_2.INIT_RAM_14 = 256'hFFFFFFC0000000000000000003FFFFFFFFFFFFE0000000000000000007FFFFFF;
defparam prom_inst_2.INIT_RAM_15 = 256'hFFFFFF80000000000000000001FFFFFFFFFFFF80000000000000000001FFFFFF;
defparam prom_inst_2.INIT_RAM_16 = 256'hFFFFFF00000000000000000000FFFFFFFFFFFF00000000000000000000FFFFFF;
defparam prom_inst_2.INIT_RAM_17 = 256'hFFFFFE000000000000000000007FFFFFFFFFFE000000000000000000007FFFFF;
defparam prom_inst_2.INIT_RAM_18 = 256'hFFFFFC000000000000000000003FFFFFFFFFFC000000000000000000003FFFFF;
defparam prom_inst_2.INIT_RAM_19 = 256'hFFFFF8000000000000000000001FFFFFFFFFFC000000000000000000003FFFFF;
defparam prom_inst_2.INIT_RAM_1A = 256'hFFFFF8000000000000000000001FFFFFFFFFF8000000000000000000001FFFFF;
defparam prom_inst_2.INIT_RAM_1B = 256'hFFFFF0000000000000000000000FFFFFFFFFF8000000000000000000001FFFFF;
defparam prom_inst_2.INIT_RAM_1C = 256'hFFFFF0000000000000000000000FFFFFFFFFF0000000000000000000000FFFFF;
defparam prom_inst_2.INIT_RAM_1D = 256'hFFFFF0000000000000000000000FFFFFFFFFF0000000000000000000000FFFFF;
defparam prom_inst_2.INIT_RAM_1E = 256'hFFFFF0000000000000000000000FFFFFFFFFF0000000000000000000000FFFFF;
defparam prom_inst_2.INIT_RAM_1F = 256'hFFFFF0000000000000000000000FFFFFFFFFF0000000000000000000000FFFFF;
defparam prom_inst_2.INIT_RAM_20 = 256'hFFFFF0000000000000000000000FFFFFFFFFF0000000000000000000000FFFFF;
defparam prom_inst_2.INIT_RAM_21 = 256'hFFFFF0000000000000000000000FFFFFFFFFF0000000000000000000000FFFFF;
defparam prom_inst_2.INIT_RAM_22 = 256'hFFFFF0000000000000000000000FFFFFFFFFF0000000000000000000000FFFFF;
defparam prom_inst_2.INIT_RAM_23 = 256'hFFFFF0000000000000000000000FFFFFFFFFF0000000000000000000000FFFFF;
defparam prom_inst_2.INIT_RAM_24 = 256'hFFFFF0000000000000000000000FFFFFFFFFF0000000000000000000000FFFFF;
defparam prom_inst_2.INIT_RAM_25 = 256'hFFFFF8000000000000000000001FFFFFFFFFF8000000000000000000001FFFFF;
defparam prom_inst_2.INIT_RAM_26 = 256'hFFFFFC000000000000000000003FFFFFFFFFF8000000000000000000001FFFFF;
defparam prom_inst_2.INIT_RAM_27 = 256'hFFFFFC000000000000000000003FFFFFFFFFFC000000000000000000003FFFFF;
defparam prom_inst_2.INIT_RAM_28 = 256'hFFFFFE000000000000000000007FFFFFFFFFFE000000000000000000007FFFFF;
defparam prom_inst_2.INIT_RAM_29 = 256'hFFFFFF00000000000000000000FFFFFFFFFFFE000000000000000000007FFFFF;
defparam prom_inst_2.INIT_RAM_2A = 256'hFFFFFF80000000000000000001FFFFFFFFFFFF00000000000000000000FFFFFF;
defparam prom_inst_2.INIT_RAM_2B = 256'hFFFFFFC0000000000000000003FFFFFFFFFFFFC0000000000000000003FFFFFF;
defparam prom_inst_2.INIT_RAM_2C = 256'hFFFFFFF000000000000000000FFFFFFFFFFFFFE0000000000000000007FFFFFF;
defparam prom_inst_2.INIT_RAM_2D = 256'hFFFFFFF800000000000000001FFFFFFFFFFFFFF000000000000000000FFFFFFF;
defparam prom_inst_2.INIT_RAM_2E = 256'hFFFFFFFE00000000000000007FFFFFFFFFFFFFFC00000000000000003FFFFFFF;
defparam prom_inst_2.INIT_RAM_2F = 256'hFFFFFFFF8000000000000001FFFFFFFFFFFFFFFF0000000000000000FFFFFFFF;
defparam prom_inst_2.INIT_RAM_30 = 256'hFFFFFFFFE000000000000007FFFFFFFFFFFFFFFFC000000000000003FFFFFFFF;
defparam prom_inst_2.INIT_RAM_31 = 256'hFFFFFFFFF80000000000001FFFFFFFFFFFFFFFFFF00000000000000FFFFFFFFF;
defparam prom_inst_2.INIT_RAM_32 = 256'hFFFFFFFFFF000000000000FFFFFFFFFFFFFFFFFFFC0000000000003FFFFFFFFF;
defparam prom_inst_2.INIT_RAM_33 = 256'hFFFFFFFFFFE00000000007FFFFFFFFFFFFFFFFFFFF800000000001FFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_34 = 256'hFFFFFFFFFFFF00000000FFFFFFFFFFFFFFFFFFFFFFF8000000001FFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_35 = 256'hFFFFFFFFFFFFFC00003FFFFFFFFFFFFFFFFFFFFFFFFFE0000007FFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00FFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[30:0],prom_inst_3_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 1;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_03 = 256'hFFFFFFFFFFFC3803FE1FFFFFFFFFFFFFFFFFFFFFFFFE003FFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_04 = 256'hFFFFFFFFFFF9FFFC01E0FFFFFFFFFFFFFFFFFFFFFFF9FFC00003FFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_05 = 256'hFFFFFFFFFFFCFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFF9FFFFFFF87FFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_06 = 256'hFFFFFFFFFFFE1FFFFFFFC7FFFFFFFFFFFFFFFFFFFFFC7FFFFFFF8FFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_07 = 256'hFFFFFFFFFFFF81E1FFFFF0FFFFFFFFFFFFFFFFFFFFFF8FFFFFFFE3FFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_08 = 256'hFFFFFFFFFFC07E0E7FFFFE3FFFFFFFFFFFFFFFFFFFF80000FFFFFC7FFFFFFFFF;
defparam prom_inst_3.INIT_RAM_09 = 256'hFFFFFFFFF03FFFCF0F1FFF8FFFFFFFFFFFFFFFFFFC07FFCF3FBFFF1FFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0A = 256'hFFFFFFFE0FFFFF87CFCFFFF3FFFFFFFFFFFFFFFF83FFFF8F801FFFE7FFFFFFFF;
defparam prom_inst_3.INIT_RAM_0B = 256'hFFFFFFF9FFFFFFB383E7FFFCFFFFFFFFFFFFFFFC7FFFFF83C7CFFFF9FFFFFFFF;
defparam prom_inst_3.INIT_RAM_0C = 256'hFFFFFFF3FFFF9F9C7C71FFFE3FFFFFFFFFFFFFF3FFFFFFB818F3FFFE7FFFFFFF;
defparam prom_inst_3.INIT_RAM_0D = 256'hFFFFFFFC3FF8439FFF3C67FF9FFFFFFFFFFFFFF8FFFE0F9FFE78E7FF3FFFFFFF;
defparam prom_inst_3.INIT_RAM_0E = 256'hFFFFFFFFC003C00FFFCF8FFFCFFFFFFFFFFFFFFE0000E00FFF9E0FFFCFFFFFFF;
defparam prom_inst_3.INIT_RAM_0F = 256'hFFFFFFFFFFF87FE7FFE79FFFE7FFFFFFFFFFFFFFFFFE0FC7FFC79FFFE7FFFFFF;
defparam prom_inst_3.INIT_RAM_10 = 256'hFFFFFFFFFF0FFFF9FFF39FFFF3FFFFFFFFFFFFFFFFC1FFF3FFF39FFFF3FFFFFF;
defparam prom_inst_3.INIT_RAM_11 = 256'hFFFFFFFFE0FFFFFE7FF9CFFFF9FFFFFFFFFFFFFFF83FFFF8FFF9CFFFFBFFFFFF;
defparam prom_inst_3.INIT_RAM_12 = 256'hFFFFFFFF1FFFFFF98FFCE7FFF9FFFFFFFFFFFFFF87FFFFFF1FFCCFFFF9FFFFFF;
defparam prom_inst_3.INIT_RAM_13 = 256'hFFFFFFFE7FFFC003CFFE73FFF9FFFFFFFFFFFFFE3FFFFFC1CFFE63FFF9FFFFFF;
defparam prom_inst_3.INIT_RAM_14 = 256'hFFFFFFFE7FFE3FFC4FFF3C3FFCFFFFFFFFFFFFFE7FFF8039EFFF399FFCFFFFFF;
defparam prom_inst_3.INIT_RAM_15 = 256'hFFFFFFFF3FE1FFFFC7FF80FFFCFFFFFFFFFFFFFE7FF87FFE07FF987FFCFFFFFF;
defparam prom_inst_3.INIT_RAM_16 = 256'hFFFFFFFF801FFFFE67FFE7FFFE7FFFFFFFFFFFFF8003FFFFE7FFC7FFFCFFFFFF;
defparam prom_inst_3.INIT_RAM_17 = 256'hFFFFFFFF9FFF7C7CF3FFF9FFFE7FFFFFFFFFFFFF9FFFFE3CF3FFF3FFFE7FFFFF;
defparam prom_inst_3.INIT_RAM_18 = 256'hFFFFFFFF9FFE00F9F1FFFE3FFF7FFFFFFFFFFFFF9FFF20FDF3FFFCFFFE7FFFFF;
defparam prom_inst_3.INIT_RAM_19 = 256'hFFFFFFFFC7F0FF09F9FFFFDFFF3FFFFFFFFFFFFF8FFC3E39F9FFFF1FFF3FFFFF;
defparam prom_inst_3.INIT_RAM_1A = 256'hFFFFFFFFF80FFFF9FCFFFFFFFF3FFFFFFFFFFFFFE001FF81FCFFFFFFFF3FFFFF;
defparam prom_inst_3.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFCFE7FFFFFFFBFFFFFFFFFFFFFFFFFFFF9FE7FFFFFFF3FFFFF;
defparam prom_inst_3.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFCCFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFCDF3FFFFFFF9FFFFF;
defparam prom_inst_3.INIT_RAM_1D = 256'hFFFFFFF807FFFFFE1FFFFFFFFF9FFFFFFFFFFFFC3FFFFFFE1FFFFFFFFF9FFFFF;
defparam prom_inst_3.INIT_RAM_1E = 256'hFFFFFFF8E01FFFFF9FFFFFFFFF9FFFFFFFFFFFF880FFFFFF1FFFFFFFFF9FFFFF;
defparam prom_inst_3.INIT_RAM_1F = 256'hF0000000FF80FFFF9FFFFFFFFFDFFFFFF0000000FC07FFFF9FFFFFFFFFDFFFFF;
defparam prom_inst_3.INIT_RAM_20 = 256'hF3FFFFFFFFFE03FF9FFFFFFFFFCFFFFFF3FFFFFFFFF01FFF9FFFFFFFFFCFFFFF;
defparam prom_inst_3.INIT_RAM_21 = 256'hF3FFFFFFFFFFF03F9FFFFFFFFFCFFFFFF3FFFFFFFFFFC07F9FFFFFFFFFCFFFFF;
defparam prom_inst_3.INIT_RAM_22 = 256'hF3FFFFFFFFFF01FF9FFFFFFFFFCFFFFFF3FFFFFFFFFFE07F9FFFFFFFFFCFFFFF;
defparam prom_inst_3.INIT_RAM_23 = 256'hF0000000FFC07FFFDFFFFFFFFFCFFFFFF3FFFFFFFFF80FFF9FFFFFFFFFCFFFFF;
defparam prom_inst_3.INIT_RAM_24 = 256'hFFFFFFF8F81FFFFFCFFFFFFFFFCFFFFFF0000000FE03FFFFCFFFFFFFFFCFFFFF;
defparam prom_inst_3.INIT_RAM_25 = 256'hFFFFFFF803FFFFFFEFFFFFFFFFCFFFFFFFFFFFF8C0FFFFFFCFFFFFFFFFCFFFFF;
defparam prom_inst_3.INIT_RAM_26 = 256'hFFFFFFFCFFFFFFFFE7FFFFFFFFCFFFFFFFFFFFF81FFFFFFFE7FFFFFFFFCFFFFF;
defparam prom_inst_3.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFF3FFFFFFFFCFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFCFFFFF;
defparam prom_inst_3.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFF9FFFFFFFFCFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFCFFFFF;
defparam prom_inst_3.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFCFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFF9FFFFFFFFCFFFFF;
defparam prom_inst_3.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFE7FFFFFFFE7FFFFFFFFFFFFFFFFFFFFFCFFFFFFFFE7FFFF;
defparam prom_inst_3.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFF3FFFFFFFF3FFFFFFFFFFFFFFFFFFFFFE7FFFFFFFF3FFFF;
defparam prom_inst_3.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFF9FFFFFFFF8FFFFFFFFFFFFFFFFFFFFFF3FFFFFFFF9FFFF;
defparam prom_inst_3.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFCFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFF9FFFFFFFFCFFFF;
defparam prom_inst_3.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFE7FFFFFFFF1FFFFFFFFFFFFFFFFFFFFFC7FFFFFFFE3FFF;
defparam prom_inst_3.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFF1FFFFFFFFC7FFFFFFFFFFFFFFFFFFFFF3FFFFFFFF8FFF;
defparam prom_inst_3.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFC7FFFFFFFF9FFFFFFFFFFFFFFFFFFFFF8FFFFFFFFE3FF;
defparam prom_inst_3.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFF1FFFFFFFFE3FFFFFFFFFFFFFFFFFFFFE3FFFFFFFFC7F;
defparam prom_inst_3.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFF3F;
defparam prom_inst_3.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0FFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFF;
defparam prom_inst_3.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFF;
defparam prom_inst_3.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFF;
defparam prom_inst_3.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFF;
defparam prom_inst_3.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFF;
defparam prom_inst_3.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFF;
defparam prom_inst_3.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[30:0],prom_inst_4_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_4),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_4.READ_MODE = 1'b0;
defparam prom_inst_4.BIT_WIDTH = 1;
defparam prom_inst_4.RESET_MODE = "SYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_03 = 256'hFFFFFFFFFFFC3807FE1FFFFFFFFFFFFFFFFFFFFFFFFE003FFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_04 = 256'hFFFFFFFFFFF9FFFC01E0FFFFFFFFFFFFFFFFFFFFFFF9FFC00003FFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_05 = 256'hFFFFFFFFFFFCFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFF9FFFFFFF87FFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_06 = 256'hFFFFFFFFFFFE1FFFFFFFC7FFFFFFFFFFFFFFFFFFFFFC7FFFFFFF8FFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_07 = 256'hFFFFFFFFFFFF81E1FFFFF0FFFFFFFFFFFFFFFFFFFFFF8FFFFFFFE3FFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_08 = 256'hFFFFFFFFFFC07E0E7FFFFE3FFFFFFFFFFFFFFFFFFFF80000FFFFFC7FFFFFFFFF;
defparam prom_inst_4.INIT_RAM_09 = 256'hFFFFFFFFF03FFFCF0F1FFF8FFFFFFFFFFFFFFFFFFC07FFCF3FBFFF1FFFFFFFFF;
defparam prom_inst_4.INIT_RAM_0A = 256'hFFFFFFFE0FFFFF87CFCFFFF3FFFFFFFFFFFFFFFF83FFFF8F801FFFE7FFFFFFFF;
defparam prom_inst_4.INIT_RAM_0B = 256'hFFFFFFF9FFFFFFB383E7FFFCFFFFFFFFFFFFFFFC7FFFFF83C7CFFFF9FFFFFFFF;
defparam prom_inst_4.INIT_RAM_0C = 256'hFFFFFFF3FFFF9F9C7C71FFFE3FFFFFFFFFFFFFF3FFFFFFB818F3FFFE7FFFFFFF;
defparam prom_inst_4.INIT_RAM_0D = 256'hFFFFFFFC3FF8439FFF3C67FF9FFFFFFFFFFFFFF8FFFE0F9FFE78E7FF3FFFFFFF;
defparam prom_inst_4.INIT_RAM_0E = 256'hFFFFFFFFC003C00FFFCF8FFFCFFFFFFFFFFFFFFE0000E00FFF9E0FFFCFFFFFFF;
defparam prom_inst_4.INIT_RAM_0F = 256'hFFFFFFFFFFF87FE7FFE79FFFE7FFFFFFFFFFFFFFFFFE0FC7FFC79FFFE7FFFFFF;
defparam prom_inst_4.INIT_RAM_10 = 256'hFFFFFFFFFF0FFFF9FFF39FFFF3FFFFFFFFFFFFFFFFC1FFF3FFF39FFFF3FFFFFF;
defparam prom_inst_4.INIT_RAM_11 = 256'hFFFFFFFFE0FFFFFE7FF9CFFFF9FFFFFFFFFFFFFFF83FFFF8FFF9CFFFFBFFFFFF;
defparam prom_inst_4.INIT_RAM_12 = 256'hFFFFFFFF1FFFFFF98FFCE7FFF9FFFFFFFFFFFFFF87FFFFFF1FFCCFFFF9FFFFFF;
defparam prom_inst_4.INIT_RAM_13 = 256'hFFFFFFFE7FFFC003CFFE73FFF9FFFFFFFFFFFFFE3FFFFFC1CFFE63FFF9FFFFFF;
defparam prom_inst_4.INIT_RAM_14 = 256'hFFFFFFFE7FFE3FFC4FFF3C3FFCFFFFFFFFFFFFFE7FFF8039EFFF399FFCFFFFFF;
defparam prom_inst_4.INIT_RAM_15 = 256'hFFFFFFFF3FE1FFFFC7FF80FFFCFFFFFFFFFFFFFE7FF87FFE07FF987FFCFFFFFF;
defparam prom_inst_4.INIT_RAM_16 = 256'hFFFFFFFF801FFFFE67FFE7FFFE7FFFFFFFFFFFFF8003FFFFE7FFC7FFFCFFFFFF;
defparam prom_inst_4.INIT_RAM_17 = 256'hFFFFFFFF9FFF7C7CF3FFF9FFFE7FFFFFFFFFFFFF9FFFFE3CF3FFF3FFFE7FFFFF;
defparam prom_inst_4.INIT_RAM_18 = 256'hFFFFFFFF9FFE00F9F1FFFE3FFF7FFFFFFFFFFFFF9FFF20FDF3FFFCFFFE7FFFFF;
defparam prom_inst_4.INIT_RAM_19 = 256'hFFFFFFFFC7F0FF09F9FFFFDFFF3FFFFFFFFFFFFF8FFC3E39F9FFFF1FFF3FFFFF;
defparam prom_inst_4.INIT_RAM_1A = 256'hFFFFFFFFF80FFFF9FCFFFFFFFF3FFFFFFFFFFFFFE001FF81FCFFFFFFFF3FFFFF;
defparam prom_inst_4.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFCFE7FFFFFFFBFFFFFFFFFFFFFFFFFFFF9FE7FFFFFFF3FFFFF;
defparam prom_inst_4.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFCCFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFCDF3FFFFFFF9FFFFF;
defparam prom_inst_4.INIT_RAM_1D = 256'hFFFFFFC07FFFFFFE1FFFFFFFFF9FFFFFFFFFFFF8FFFFFFFE1FFFFFFFFF9FFFFF;
defparam prom_inst_4.INIT_RAM_1E = 256'hFFFFF80C7FFFFFFF9FFFFFFFFF9FFFFFFFFFFF007FFFFFFF1FFFFFFFFF9FFFFF;
defparam prom_inst_4.INIT_RAM_1F = 256'hFFFE03FC0000003F9FFFFFFFFFDFFFFFFFFFC07C7FFFFFFF9FFFFFFFFFDFFFFF;
defparam prom_inst_4.INIT_RAM_20 = 256'hFF80FFFFFFFFFF3F9FFFFFFFFFCFFFFFFFF01FFE0000003F9FFFFFFFFFCFFFFF;
defparam prom_inst_4.INIT_RAM_21 = 256'hF01FFFFFFFFFFF3F9FFFFFFFFFCFFFFFFC03FFFFFFFFFF3F9FFFFFFFFFCFFFFF;
defparam prom_inst_4.INIT_RAM_22 = 256'hF80FFFFFFFFFFF3F9FFFFFFFFFCFFFFFF03FFFFFFFFFFF3F9FFFFFFFFFCFFFFF;
defparam prom_inst_4.INIT_RAM_23 = 256'hFFF03FFE0000003FDFFFFFFFFFCFFFFFFF81FFFFFFFFFF3F9FFFFFFFFFCFFFFF;
defparam prom_inst_4.INIT_RAM_24 = 256'hFFFF80FC0000003FCFFFFFFFFFCFFFFFFFFC07FC0000003FCFFFFFFFFFCFFFFF;
defparam prom_inst_4.INIT_RAM_25 = 256'hFFFFFE007FFFFFFFEFFFFFFFFFCFFFFFFFFFF01C7FFFFFFFCFFFFFFFFFCFFFFF;
defparam prom_inst_4.INIT_RAM_26 = 256'hFFFFFFF8FFFFFFFFE7FFFFFFFFCFFFFFFFFFFFC07FFFFFFFE7FFFFFFFFCFFFFF;
defparam prom_inst_4.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFF3FFFFFFFFCFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFCFFFFF;
defparam prom_inst_4.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFF9FFFFFFFFCFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFCFFFFF;
defparam prom_inst_4.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFCFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFF9FFFFFFFFCFFFFF;
defparam prom_inst_4.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFE7FFFFFFFE7FFFFFFFFFFFFFFFFFFFFFCFFFFFFFFE7FFFF;
defparam prom_inst_4.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFF3FFFFFFFF3FFFFFFFFFFFFFFFFFFFFFE7FFFFFFFF3FFFF;
defparam prom_inst_4.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFF9FFFFFFFF8FFFFFFFFFFFFFFFFFFFFFF3FFFFFFFF9FFFF;
defparam prom_inst_4.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFCFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFF9FFFFFFFFCFFFF;
defparam prom_inst_4.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFE7FFFFFFFF1FFFFFFFFFFFFFFFFFFFFFC7FFFFFFFE3FFF;
defparam prom_inst_4.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFF1FFFFFFFFC7FFFFFFFFFFFFFFFFFFFFF3FFFFFFFF8FFF;
defparam prom_inst_4.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFC7FFFFFFFF9FFFFFFFFFFFFFFFFFFFFF8FFFFFFFFE3FF;
defparam prom_inst_4.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFF1FFFFFFFFE3FFFFFFFFFFFFFFFFFFFFE3FFFFFFFFC7F;
defparam prom_inst_4.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFF3F;
defparam prom_inst_4.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0FFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFF;
defparam prom_inst_4.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFF;
defparam prom_inst_4.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFF;
defparam prom_inst_4.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFF;
defparam prom_inst_4.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFF;
defparam prom_inst_4.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFF;
defparam prom_inst_4.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[30:0],prom_inst_5_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_5),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_5.READ_MODE = 1'b0;
defparam prom_inst_5.BIT_WIDTH = 1;
defparam prom_inst_5.RESET_MODE = "SYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_08 = 256'hFFFFFFFFFFFFF000000FFFFFFFFFFFFFFFFFFFFFFFFFFFE007FFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_09 = 256'hFFFFFFFFFFF8000000001FFFFFFFFFFFFFFFFFFFFFFF00000000FFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_0A = 256'hFFFFFFFFFF000FFFFFF001FFFFFFFFFFFFFFFFFFFFE0003FFC0007FFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_0B = 256'hFFFFFFFFF003FFFFFFFFC01FFFFFFFFFFFFFFFFFFC00FFFFFFFE003FFFFFFFFF;
defparam prom_inst_5.INIT_RAM_0C = 256'hFFFFFFFF807FFFFFFFFFFE01FFFFFFFFFFFFFFFFE01FFFFFFFFFF807FFFFFFFF;
defparam prom_inst_5.INIT_RAM_0D = 256'hFFFFFFFE07FFFFFFFFFFFFC07FFFFFFFFFFFFFFF01FFFFFFFFFFFF80FFFFFFFF;
defparam prom_inst_5.INIT_RAM_0E = 256'hFFFFFFF03FFFFFF00FFFFFF80FFFFFFFFFFFFFF80FFFFFFFFFFFFFF01FFFFFFF;
defparam prom_inst_5.INIT_RAM_0F = 256'hFFFFFFC0FFFFE0000007FFFF03FFFFFFFFFFFFE07FFFFC00003FFFFE07FFFFFF;
defparam prom_inst_5.INIT_RAM_10 = 256'hFFFFFF03FFFC000000003FFFC0FFFFFFFFFFFF81FFFF00000000FFFF81FFFFFF;
defparam prom_inst_5.INIT_RAM_11 = 256'hFFFFFC1FFFC00000000003FFF03FFFFFFFFFFE0FFFF0000000000FFFE07FFFFF;
defparam prom_inst_5.INIT_RAM_12 = 256'hFFFFF83FFE0000000000007FFC1FFFFFFFFFF81FFF800000000001FFF81FFFFF;
defparam prom_inst_5.INIT_RAM_13 = 256'hFFFFE0FFF80000000000001FFF07FFFFFFFFF07FFC0000000000003FFE0FFFFF;
defparam prom_inst_5.INIT_RAM_14 = 256'hFFFFC1FFE000000000000007FF83FFFFFFFFC1FFF00000000000000FFF87FFFF;
defparam prom_inst_5.INIT_RAM_15 = 256'hFFFF87FF8003F000000F8001FFE1FFFFFFFF83FFC001E00000070003FFC1FFFF;
defparam prom_inst_5.INIT_RAM_16 = 256'hFFFF0FFE0003FC00003FC0007FF0FFFFFFFF07FF0003F800001FC000FFE0FFFF;
defparam prom_inst_5.INIT_RAM_17 = 256'hFFFE1FFC0001FF0000FF80003FF87FFFFFFE0FFE0003FE00007FC0007FF07FFF;
defparam prom_inst_5.INIT_RAM_18 = 256'hFFFC3FF800007FC003FE00001FFC3FFFFFFC1FF80000FF8001FF00001FF83FFF;
defparam prom_inst_5.INIT_RAM_19 = 256'hFFF87FF000001FF00FF800000FFE1FFFFFF83FF000003FE007FC00000FFC3FFF;
defparam prom_inst_5.INIT_RAM_1A = 256'hFFF07FE0000007FC3FE0000007FE1FFFFFF87FE000000FF81FF0000007FE1FFF;
defparam prom_inst_5.INIT_RAM_1B = 256'hFFF0FFC0000001FFFF80000003FF0FFFFFF0FFC0000003FE7FC0000003FF0FFF;
defparam prom_inst_5.INIT_RAM_1C = 256'hFFE1FF800000007FFE00000001FF07FFFFF0FFC0000000FFFF00000003FF0FFF;
defparam prom_inst_5.INIT_RAM_1D = 256'hFFE1FF800000FFFFFFFF000001FF87FFFFE1FF800000003FFC00000001FF87FF;
defparam prom_inst_5.INIT_RAM_1E = 256'hFFE1FF000003FFFFFFFFC00000FF87FFFFE1FF800001FFFFFFFF800001FF87FF;
defparam prom_inst_5.INIT_RAM_1F = 256'hFFC3FF000003FFFFFFFFC00000FF87FFFFE1FF000003FFFFFFFFC00000FF87FF;
defparam prom_inst_5.INIT_RAM_20 = 256'hFFC3FF0000007FFFFFFE000000FFC3FFFFC3FF000001FFFFFFFF800000FF83FF;
defparam prom_inst_5.INIT_RAM_21 = 256'hFFC3FF0000000007E000000000FFC3FFFFC3FF0000000007E000000000FFC3FF;
defparam prom_inst_5.INIT_RAM_22 = 256'hFFC3FF0000000007E000000000FFC3FFFFC3FF0000000007E000000000FFC3FF;
defparam prom_inst_5.INIT_RAM_23 = 256'hFFC3FF000001FFFFFFFF800000FFC3FFFFC3FF0000000007E000000000FFC3FF;
defparam prom_inst_5.INIT_RAM_24 = 256'hFFC1FF000003FFFFFFFFC00000FF87FFFFC3FF000003FFFFFFFFC00000FF87FF;
defparam prom_inst_5.INIT_RAM_25 = 256'hFFE1FF000003FFFFFFFF800001FF87FFFFE1FF000003FFFFFFFFC00000FF87FF;
defparam prom_inst_5.INIT_RAM_26 = 256'hFFE1FF8000000007E000000001FF87FFFFE1FF800001FFFFFFFF000001FF87FF;
defparam prom_inst_5.INIT_RAM_27 = 256'hFFF0FFC000000007E000000003FF0FFFFFE1FF8000000007E000000001FF07FF;
defparam prom_inst_5.INIT_RAM_28 = 256'hFFF0FFC000000007E000000003FF0FFFFFF0FFC000000007E000000003FF0FFF;
defparam prom_inst_5.INIT_RAM_29 = 256'hFFF87FE000000007E000000007FE1FFFFFF07FE000000007E000000007FE0FFF;
defparam prom_inst_5.INIT_RAM_2A = 256'hFFF83FF000000007E00000000FFC1FFFFFF87FE000000007E00000000FFE1FFF;
defparam prom_inst_5.INIT_RAM_2B = 256'hFFFC3FF800000007E00000001FF83FFFFFFC3FF800000007E00000001FFC3FFF;
defparam prom_inst_5.INIT_RAM_2C = 256'hFFFE1FFC00000007E00000007FF07FFFFFFC1FFC00000007E00000003FF87FFF;
defparam prom_inst_5.INIT_RAM_2D = 256'hFFFF07FF00000007E0000000FFE0FFFFFFFE0FFE00000007E00000007FF0FFFF;
defparam prom_inst_5.INIT_RAM_2E = 256'hFFFF83FFC0000003C0000003FFC1FFFFFFFF07FF80000007E0000001FFE1FFFF;
defparam prom_inst_5.INIT_RAM_2F = 256'hFFFFC1FFE00000000000000FFF83FFFFFFFFC3FFC000000000000007FF83FFFF;
defparam prom_inst_5.INIT_RAM_30 = 256'hFFFFF07FFC0000000000003FFE0FFFFFFFFFE0FFF80000000000001FFF07FFFF;
defparam prom_inst_5.INIT_RAM_31 = 256'hFFFFF83FFF000000000000FFFC1FFFFFFFFFF07FFE0000000000007FFC1FFFFF;
defparam prom_inst_5.INIT_RAM_32 = 256'hFFFFFE0FFFE0000000000FFFF07FFFFFFFFFFC1FFFC00000000003FFF83FFFFF;
defparam prom_inst_5.INIT_RAM_33 = 256'hFFFFFF800FFE00000000FFFF81FFFFFFFFFFFF003FF8000000001FFFE0FFFFFF;
defparam prom_inst_5.INIT_RAM_34 = 256'hFFFFFFC003FFF800003FFFFE07FFFFFFFFFFFFC007FFC0000003FFFF03FFFFFF;
defparam prom_inst_5.INIT_RAM_35 = 256'hFFFFFF8003FFFFFFFFFFFFF01FFFFFFFFFFFFF8003FFFFC003FFFFFC0FFFFFFF;
defparam prom_inst_5.INIT_RAM_36 = 256'hFFFFFF8003FFFFFFFFFFFF80FFFFFFFFFFFFFF8001FFFFFFFFFFFFE03FFFFFFF;
defparam prom_inst_5.INIT_RAM_37 = 256'hFFFFFFC003FFFFFFFFFFF807FFFFFFFFFFFFFF8003FFFFFFFFFFFE01FFFFFFFF;
defparam prom_inst_5.INIT_RAM_38 = 256'hFFFFFFF00FFFFFFFFFFF003FFFFFFFFFFFFFFFE007FFFFFFFFFFE00FFFFFFFFF;
defparam prom_inst_5.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFF0003FFFFFFFFFFFFFFFFF83FFFFFFFFFF800FFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFF80000FFFFFFFFFFFFFFFFFFFFFFFFFFFC00001FFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_6 (
    .DO({prom_inst_6_dout_w[30:0],prom_inst_6_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_6),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_6.READ_MODE = 1'b0;
defparam prom_inst_6.BIT_WIDTH = 1;
defparam prom_inst_6.RESET_MODE = "SYNC";
defparam prom_inst_6.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFF03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF87FFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE01FFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_04 = 256'hFFFFFFFFFFFFFF800FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00FFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_05 = 256'hFFFFFFFFFFFFFF8007FFFFFFFFFFFFFFFFFFFFFFFFFFFF8007FFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_06 = 256'hFFFFFFFFFFFFFF0003FFFFFFFFFFFFFFFFFFFFFFFFFFFF0003FFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_07 = 256'hFFFFFFFFFFFFFE0301FFFFFFFFFFFFFFFFFFFFFFFFFFFE0301FFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_08 = 256'hFFFFFFFFFFFFFC0780FFFFFFFFFFFFFFFFFFFFFFFFFFFC0700FFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_09 = 256'hFFFFFFFFFFFFF80FC07FFFFFFFFFFFFFFFFFFFFFFFFFF80F80FFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_0A = 256'hFFFFFFFFFFFFF01FE03FFFFFFFFFFFFFFFFFFFFFFFFFF01FC07FFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_0B = 256'hFFFFFFFFFFFFE03FF01FFFFFFFFFFFFFFFFFFFFFFFFFF01FE03FFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_0C = 256'hFFFFFFFFFFFFC07FF80FFFFFFFFFFFFFFFFFFFFFFFFFE03FF01FFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_0D = 256'hFFFFFFFFFFFF80FFF807FFFFFFFFFFFFFFFFFFFFFFFFC07FF80FFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_0E = 256'hFFFFFFFFFFFF01FFFC07FFFFFFFFFFFFFFFFFFFFFFFF80FFFC07FFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_0F = 256'hFFFFFFFFFFFE03FFFE03FFFFFFFFFFFFFFFFFFFFFFFF01FFFE03FFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_10 = 256'hFFFFFFFFFFFE03FFFF01FFFFFFFFFFFFFFFFFFFFFFFE03FFFF01FFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_11 = 256'hFFFFFFFFFFFC07FFFF80FFFFFFFFFFFFFFFFFFFFFFFC07FFFF80FFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_12 = 256'hFFFFFFFFFFF80FF01FC07FFFFFFFFFFFFFFFFFFFFFF80FF83FC07FFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_13 = 256'hFFFFFFFFFFF01FE00FE03FFFFFFFFFFFFFFFFFFFFFF01FE01FE03FFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_14 = 256'hFFFFFFFFFFE03FC00FF01FFFFFFFFFFFFFFFFFFFFFE03FE00FE03FFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_15 = 256'hFFFFFFFFFFC07FC00FF80FFFFFFFFFFFFFFFFFFFFFC07FC00FF01FFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_16 = 256'hFFFFFFFFFF80FFC00FFC07FFFFFFFFFFFFFFFFFFFF807FC00FF80FFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_17 = 256'hFFFFFFFFFF01FFE00FFE03FFFFFFFFFFFFFFFFFFFF80FFC00FFC07FFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_18 = 256'hFFFFFFFFFE03FFE00FFF01FFFFFFFFFFFFFFFFFFFF01FFE00FFE03FFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_19 = 256'hFFFFFFFFFC07FFE00FFF01FFFFFFFFFFFFFFFFFFFE03FFE00FFF01FFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1A = 256'hFFFFFFFFF80FFFE01FFF80FFFFFFFFFFFFFFFFFFFC07FFE01FFF80FFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1B = 256'hFFFFFFFFF00FFFF01FFFC07FFFFFFFFFFFFFFFFFF80FFFE01FFFC07FFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1C = 256'hFFFFFFFFF01FFFF01FFFE03FFFFFFFFFFFFFFFFFF01FFFF01FFFE03FFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1D = 256'hFFFFFFFFE03FFFF01FFFF01FFFFFFFFFFFFFFFFFE03FFFF01FFFF01FFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1E = 256'hFFFFFFFFC07FFFF03FFFF80FFFFFFFFFFFFFFFFFC07FFFF03FFFF80FFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1F = 256'hFFFFFFFF80FFFFF83FFFFC07FFFFFFFFFFFFFFFF80FFFFF83FFFF80FFFFFFFFF;
defparam prom_inst_6.INIT_RAM_20 = 256'hFFFFFFFF01FFFFF83FFFFE03FFFFFFFFFFFFFFFF01FFFFF83FFFFC07FFFFFFFF;
defparam prom_inst_6.INIT_RAM_21 = 256'hFFFFFFFE03FFFFF83FFFFF01FFFFFFFFFFFFFFFE01FFFFF83FFFFE03FFFFFFFF;
defparam prom_inst_6.INIT_RAM_22 = 256'hFFFFFFFC07FFFFF87FFFFF80FFFFFFFFFFFFFFFE03FFFFF87FFFFF01FFFFFFFF;
defparam prom_inst_6.INIT_RAM_23 = 256'hFFFFFFF80FFFFFF87FFFFFC07FFFFFFFFFFFFFFC07FFFFF87FFFFF80FFFFFFFF;
defparam prom_inst_6.INIT_RAM_24 = 256'hFFFFFFF01FFFFFFC7FFFFFC07FFFFFFFFFFFFFF80FFFFFF87FFFFFC07FFFFFFF;
defparam prom_inst_6.INIT_RAM_25 = 256'hFFFFFFE03FFFFFFC7FFFFFE03FFFFFFFFFFFFFF01FFFFFFC7FFFFFE03FFFFFFF;
defparam prom_inst_6.INIT_RAM_26 = 256'hFFFFFFC07FFFFFFCFFFFFFF01FFFFFFFFFFFFFE03FFFFFFCFFFFFFF01FFFFFFF;
defparam prom_inst_6.INIT_RAM_27 = 256'hFFFFFFC07FFFFFFCFFFFFFF80FFFFFFFFFFFFFC07FFFFFFCFFFFFFF80FFFFFFF;
defparam prom_inst_6.INIT_RAM_28 = 256'hFFFFFF80FFFFFFFCFFFFFFFC07FFFFFFFFFFFF80FFFFFFFCFFFFFFFC07FFFFFF;
defparam prom_inst_6.INIT_RAM_29 = 256'hFFFFFF01FFFFFFFCFFFFFFFE03FFFFFFFFFFFF01FFFFFFFCFFFFFFFE03FFFFFF;
defparam prom_inst_6.INIT_RAM_2A = 256'hFFFFFE03FFFFFFFEFFFFFFFF01FFFFFFFFFFFE03FFFFFFFEFFFFFFFE03FFFFFF;
defparam prom_inst_6.INIT_RAM_2B = 256'hFFFFFC07FFFFFFFFFFFFFFFF80FFFFFFFFFFFC07FFFFFFFEFFFFFFFF01FFFFFF;
defparam prom_inst_6.INIT_RAM_2C = 256'hFFFFF80FFFFFFFFFFFFFFFFFC07FFFFFFFFFF80FFFFFFFFFFFFFFFFF80FFFFFF;
defparam prom_inst_6.INIT_RAM_2D = 256'hFFFFF01FFFFFFFFFFFFFFFFFE03FFFFFFFFFF80FFFFFFFFFFFFFFFFFC07FFFFF;
defparam prom_inst_6.INIT_RAM_2E = 256'hFFFFE03FFFFFFFFFFFFFFFFFF01FFFFFFFFFF01FFFFFFFFFFFFFFFFFE03FFFFF;
defparam prom_inst_6.INIT_RAM_2F = 256'hFFFFC07FFFFFFFFFFFFFFFFFF00FFFFFFFFFE03FFFFFFFFFFFFFFFFFF01FFFFF;
defparam prom_inst_6.INIT_RAM_30 = 256'hFFFF80FFFFFFFFFFFFFFFFFFF80FFFFFFFFFC07FFFFFFFFFFFFFFFFFF80FFFFF;
defparam prom_inst_6.INIT_RAM_31 = 256'hFFFF01FFFFFFFFF87FFFFFFFFC07FFFFFFFF80FFFFFFFFFFFFFFFFFFFC07FFFF;
defparam prom_inst_6.INIT_RAM_32 = 256'hFFFF01FFFFFFFFE01FFFFFFFFE03FFFFFFFF01FFFFFFFFF01FFFFFFFFE03FFFF;
defparam prom_inst_6.INIT_RAM_33 = 256'hFFFE03FFFFFFFFC00FFFFFFFFF01FFFFFFFE03FFFFFFFFE00FFFFFFFFF01FFFF;
defparam prom_inst_6.INIT_RAM_34 = 256'hFFFC07FFFFFFFFC00FFFFFFFFF80FFFFFFFC07FFFFFFFFC00FFFFFFFFF80FFFF;
defparam prom_inst_6.INIT_RAM_35 = 256'hFFF80FFFFFFFFFE00FFFFFFFFFC07FFFFFF80FFFFFFFFFC00FFFFFFFFF80FFFF;
defparam prom_inst_6.INIT_RAM_36 = 256'hFFF01FFFFFFFFFF01FFFFFFFFFE03FFFFFF01FFFFFFFFFE01FFFFFFFFFC07FFF;
defparam prom_inst_6.INIT_RAM_37 = 256'hFFE03FFFFFFFFFFFFFFFFFFFFFF01FFFFFE03FFFFFFFFFF83FFFFFFFFFE03FFF;
defparam prom_inst_6.INIT_RAM_38 = 256'hFFC07FFFFFFFFFFFFFFFFFFFFFF80FFFFFE03FFFFFFFFFFFFFFFFFFFFFF01FFF;
defparam prom_inst_6.INIT_RAM_39 = 256'hFFC07FFFFFFFFFFFFFFFFFFFFFF80FFFFFC07FFFFFFFFFFFFFFFFFFFFFF80FFF;
defparam prom_inst_6.INIT_RAM_3A = 256'hFF8000000000000000000000000007FFFFC000000000000000000000000007FF;
defparam prom_inst_6.INIT_RAM_3B = 256'hFFC000000000000000000000000007FFFF8000000000000000000000000007FF;
defparam prom_inst_6.INIT_RAM_3C = 256'hFFC00000000000000000000000000FFFFFC000000000000000000000000007FF;
defparam prom_inst_6.INIT_RAM_3D = 256'hFFF00000000000000000000000003FFFFFE00000000000000000000000000FFF;
defparam prom_inst_6.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_7 (
    .DO({prom_inst_7_dout_w[30:0],prom_inst_7_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_7),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_7.READ_MODE = 1'b0;
defparam prom_inst_7.BIT_WIDTH = 1;
defparam prom_inst_7.RESET_MODE = "SYNC";
defparam prom_inst_7.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_0A = 256'hFFFFFFFFFFFFF000000FFFFFFFFFFFFFFFFFFFFFFFFFFF8001FFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_0B = 256'hFFFFFFFFFFFC000000003FFFFFFFFFFFFFFFFFFFFFFF80000001FFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_0C = 256'hFFFFFFFFFFC00000000003FFFFFFFFFFFFFFFFFFFFF0000000000FFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_0D = 256'hFFFFFFFFFE0000000000007FFFFFFFFFFFFFFFFFFF800000000001FFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_0E = 256'hFFFFFFFFF00000000000000FFFFFFFFFFFFFFFFFFC0000000000003FFFFFFFFF;
defparam prom_inst_7.INIT_RAM_0F = 256'hFFFFFFFFC000000000000003FFFFFFFFFFFFFFFFE000000000000007FFFFFFFF;
defparam prom_inst_7.INIT_RAM_10 = 256'hFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF8000000000000001FFFFFFFF;
defparam prom_inst_7.INIT_RAM_11 = 256'hFFFFFFFC00000000000000003FFFFFFFFFFFFFFE00000000000000007FFFFFFF;
defparam prom_inst_7.INIT_RAM_12 = 256'hFFFFFFF800000000000000001FFFFFFFFFFFFFF800000000000000001FFFFFFF;
defparam prom_inst_7.INIT_RAM_13 = 256'hFFFFFFE0000000000000000007FFFFFFFFFFFFF000000000000000000FFFFFFF;
defparam prom_inst_7.INIT_RAM_14 = 256'hFFFFFFC0000000000000000003FFFFFFFFFFFFE0000000000000000007FFFFFF;
defparam prom_inst_7.INIT_RAM_15 = 256'hFFFFFF80000000000000000001FFFFFFFFFFFF80000000000000000001FFFFFF;
defparam prom_inst_7.INIT_RAM_16 = 256'hFFFFFF00000000000000000000FFFFFFFFFFFF00000000000000000000FFFFFF;
defparam prom_inst_7.INIT_RAM_17 = 256'hFFFFFE000000000000000000007FFFFFFFFFFE000000000000000000007FFFFF;
defparam prom_inst_7.INIT_RAM_18 = 256'hFFFFFC000000000000000000003FFFFFFFFFFC000000000000000000003FFFFF;
defparam prom_inst_7.INIT_RAM_19 = 256'hFFFFF8000000000000000000001FFFFFFFFFFC000000000000000000003FFFFF;
defparam prom_inst_7.INIT_RAM_1A = 256'hFFFFF8000000000000000000001FFFFFFFFFF8000000000000000000001FFFFF;
defparam prom_inst_7.INIT_RAM_1B = 256'hFFFFF0000000000000000000000FFFFFFFFFF8000000000000000000001FFFFF;
defparam prom_inst_7.INIT_RAM_1C = 256'hFFFFF0000000000000000000000FFFFFFFFFF0000000000000000000000FFFFF;
defparam prom_inst_7.INIT_RAM_1D = 256'hFFFFF0000000000000000000000FFFFFFFFFF0000000000000000000000FFFFF;
defparam prom_inst_7.INIT_RAM_1E = 256'hFFFFF0000000000000000000000FFFFFFFFFF0000000000000000000000FFFFF;
defparam prom_inst_7.INIT_RAM_1F = 256'hFFFFF0000000000000000000000FFFFFFFFFF0000000000000000000000FFFFF;
defparam prom_inst_7.INIT_RAM_20 = 256'hFFFFF0000000000000000000000FFFFFFFFFF0000000000000000000000FFFFF;
defparam prom_inst_7.INIT_RAM_21 = 256'hFFFFF0000000000000000000000FFFFFFFFFF0000000000000000000000FFFFF;
defparam prom_inst_7.INIT_RAM_22 = 256'hFFFFF0000000000000000000000FFFFFFFFFF0000000000000000000000FFFFF;
defparam prom_inst_7.INIT_RAM_23 = 256'hFFFFF0000000000000000000000FFFFFFFFFF0000000000000000000000FFFFF;
defparam prom_inst_7.INIT_RAM_24 = 256'hFFFFF0000000000000000000000FFFFFFFFFF0000000000000000000000FFFFF;
defparam prom_inst_7.INIT_RAM_25 = 256'hFFFFF8000000000000000000001FFFFFFFFFF8000000000000000000001FFFFF;
defparam prom_inst_7.INIT_RAM_26 = 256'hFFFFFC000000000000000000003FFFFFFFFFF8000000000000000000001FFFFF;
defparam prom_inst_7.INIT_RAM_27 = 256'hFFFFFC000000000000000000003FFFFFFFFFFC000000000000000000003FFFFF;
defparam prom_inst_7.INIT_RAM_28 = 256'hFFFFFE000000000000000000007FFFFFFFFFFE000000000000000000007FFFFF;
defparam prom_inst_7.INIT_RAM_29 = 256'hFFFFFF00000000000000000000FFFFFFFFFFFE000000000000000000007FFFFF;
defparam prom_inst_7.INIT_RAM_2A = 256'hFFFFFF80000000000000000001FFFFFFFFFFFF00000000000000000000FFFFFF;
defparam prom_inst_7.INIT_RAM_2B = 256'hFFFFFFC0000000000000000003FFFFFFFFFFFFC0000000000000000003FFFFFF;
defparam prom_inst_7.INIT_RAM_2C = 256'hFFFFFFF000000000000000000FFFFFFFFFFFFFE0000000000000000007FFFFFF;
defparam prom_inst_7.INIT_RAM_2D = 256'hFFFFFFF800000000000000001FFFFFFFFFFFFFF000000000000000000FFFFFFF;
defparam prom_inst_7.INIT_RAM_2E = 256'hFFFFFFFE00000000000000007FFFFFFFFFFFFFFC00000000000000003FFFFFFF;
defparam prom_inst_7.INIT_RAM_2F = 256'hFFFFFFFF8000000000000001FFFFFFFFFFFFFFFF0000000000000000FFFFFFFF;
defparam prom_inst_7.INIT_RAM_30 = 256'hFFFFFFFFE000000000000007FFFFFFFFFFFFFFFFC000000000000003FFFFFFFF;
defparam prom_inst_7.INIT_RAM_31 = 256'hFFFFFFFFF80000000000001FFFFFFFFFFFFFFFFFF00000000000000FFFFFFFFF;
defparam prom_inst_7.INIT_RAM_32 = 256'hFFFFFFFFFF000000000000FFFFFFFFFFFFFFFFFFFC0000000000003FFFFFFFFF;
defparam prom_inst_7.INIT_RAM_33 = 256'hFFFFFFFFFFE00000000007FFFFFFFFFFFFFFFFFFFF800000000001FFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_34 = 256'hFFFFFFFFFFFF00000000FFFFFFFFFFFFFFFFFFFFFFF8000000001FFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_35 = 256'hFFFFFFFFFFFFFC00003FFFFFFFFFFFFFFFFFFFFFFFFFE0000007FFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00FFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[16]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(ad[15]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_1_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(prom_inst_2_dout[0]),
  .I1(prom_inst_3_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(prom_inst_4_dout[0]),
  .I1(prom_inst_5_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(prom_inst_6_dout[0]),
  .I1(prom_inst_7_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_1)
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(dff_q_1)
);
MUX2 mux_inst_6 (
  .O(dout[0]),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(dff_q_0)
);
endmodule //ROM_picture
