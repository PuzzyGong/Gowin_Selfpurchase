`include "../define.v"

module uart_sfr
(
    input  wire                         sys_clk                    ,
    input  wire                         sys_rst_n                  ,

    input  wire                         rx                         ,
    output wire                         tx                         ,
    output wire        [256-1:0]        o_contains                  
);

wire                   [   7:0]         data                       ;
wire                   [  15:0]         address                    ;
wire                                    ad_set                     ;
wire                                    ad_enable                  ;

debug u_debug(
    .sys_clk                           (sys_clk                   ),
    .sys_rst_n                         (sys_rst_n                 ),
    .data_io                           (data                      ),
    .d_address                         (address                   ),
    .d_set                             (ad_set                    ),
    .d_enable                          (ad_enable                 ),
    .rx                                (rx                        ),
    .tx                                (tx                        ) 
);

//**************************** sfr ****************************

sfr#(.RST_VALUE                         (`RST_VALUE_0000           ),                        .SFR_ADDRESS                       (16'h00                     )                         )                       u_sfr00(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h00,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_0001           ),                        .SFR_ADDRESS                       (16'h01                     )                         )                       u_sfr01(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h01,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_0002           ),                        .SFR_ADDRESS                       (16'h02                     )                         )                       u_sfr02(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h02,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_0003           ),                        .SFR_ADDRESS                       (16'h03                     )                         )                       u_sfr03(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h03,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_0004           ),                        .SFR_ADDRESS                       (16'h04                     )                         )                       u_sfr04(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h04,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_0005           ),                        .SFR_ADDRESS                       (16'h05                     )                         )                       u_sfr05(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h05,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_0006           ),                        .SFR_ADDRESS                       (16'h06                     )                         )                       u_sfr06(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h06,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_0007           ),                        .SFR_ADDRESS                       (16'h07                     )                         )                       u_sfr07(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h07,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_0008           ),                        .SFR_ADDRESS                       (16'h08                     )                         )                       u_sfr08(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h08,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_0009           ),                        .SFR_ADDRESS                       (16'h09                     )                         )                       u_sfr09(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h09,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_000A           ),                        .SFR_ADDRESS                       (16'h0A                     )                         )                       u_sfr0A(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h0A,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_000B           ),                        .SFR_ADDRESS                       (16'h0B                     )                         )                       u_sfr0B(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h0B,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_000C           ),                        .SFR_ADDRESS                       (16'h0C                     )                         )                       u_sfr0C(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h0C,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_000D           ),                        .SFR_ADDRESS                       (16'h0D                     )                         )                       u_sfr0D(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h0D,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_000E           ),                        .SFR_ADDRESS                       (16'h0E                     )                         )                       u_sfr0E(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h0E,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_000F           ),                        .SFR_ADDRESS                       (16'h0F                     )                         )                       u_sfr0F(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h0F,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_0010           ),                        .SFR_ADDRESS                       (16'h10                     )                         )                       u_sfr10(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h10,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_0011           ),                        .SFR_ADDRESS                       (16'h11                     )                         )                       u_sfr11(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h11,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_0012           ),                        .SFR_ADDRESS                       (16'h12                     )                         )                       u_sfr12(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h12,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_0013           ),                        .SFR_ADDRESS                       (16'h13                     )                         )                       u_sfr13(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h13,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_0014           ),                        .SFR_ADDRESS                       (16'h14                     )                         )                       u_sfr14(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h14,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_0015           ),                        .SFR_ADDRESS                       (16'h15                     )                         )                       u_sfr15(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h15,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_0016           ),                        .SFR_ADDRESS                       (16'h16                     )                         )                       u_sfr16(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h16,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_0017           ),                        .SFR_ADDRESS                       (16'h17                     )                         )                       u_sfr17(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h17,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_0018           ),                        .SFR_ADDRESS                       (16'h18                     )                         )                       u_sfr18(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h18,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_0019           ),                        .SFR_ADDRESS                       (16'h19                     )                         )                       u_sfr19(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h19,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_001A           ),                        .SFR_ADDRESS                       (16'h1A                     )                         )                       u_sfr1A(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h1A,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_001B           ),                        .SFR_ADDRESS                       (16'h1B                     )                         )                       u_sfr1B(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h1B,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_001C           ),                        .SFR_ADDRESS                       (16'h1C                     )                         )                       u_sfr1C(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h1C,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_001D           ),                        .SFR_ADDRESS                       (16'h1D                     )                         )                       u_sfr1D(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h1D,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_001E           ),                        .SFR_ADDRESS                       (16'h1E                     )                         )                       u_sfr1E(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h1E,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );
sfr#(.RST_VALUE                         (`RST_VALUE_001F           ),                        .SFR_ADDRESS                       (16'h1F                     )                         )                       u_sfr1F(                     .sys_clk                           (sys_clk                   ),                        .sys_rst_n                         (sys_rst_n                 ),                        .i_address                         (address                   ),                        .i_ad_set                          (ad_set                    ),                        .i_ad_enable                       (ad_enable                 ),                        .io_ad_data                        (data                      ),                        .i_set                             (1'b0                      ),                        .i_enable                          (1'b0                      ),                        .i_data                            (8'd0                      ),                        .o_data                            (                          ),                        .o_contain                         (o_contains[{'h1F,3'd0}+:8]   ),                        .o_rd_flag                         (                          ),                        .o_wt_flag                         (                          )                         );


endmodule